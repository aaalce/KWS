// This is the unpowered netlist.
module kws_wrapper (wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i);
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;

 wire net59;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire clknet_0_wb_clk_i;
 wire clknet_2_0__leaf_wb_clk_i;
 wire clknet_2_1__leaf_wb_clk_i;
 wire clknet_2_2__leaf_wb_clk_i;
 wire clknet_2_3__leaf_wb_clk_i;
 wire \fsm_inst.batch_norm_en ;
 wire \fsm_inst.cnn_en ;
 wire \fsm_inst.current_state[0] ;
 wire \fsm_inst.current_state[1] ;
 wire \fsm_inst.current_state[2] ;
 wire \fsm_inst.done ;
 wire \fsm_inst.next_state[0] ;
 wire \fsm_inst.next_state[1] ;
 wire \fsm_inst.next_state[2] ;
 wire net1;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net9;
 wire \weights_inst.data_out[0] ;
 wire \weights_inst.data_out[10] ;
 wire \weights_inst.data_out[11] ;
 wire \weights_inst.data_out[12] ;
 wire \weights_inst.data_out[13] ;
 wire \weights_inst.data_out[14] ;
 wire \weights_inst.data_out[15] ;
 wire \weights_inst.data_out[16] ;
 wire \weights_inst.data_out[17] ;
 wire \weights_inst.data_out[18] ;
 wire \weights_inst.data_out[19] ;
 wire \weights_inst.data_out[1] ;
 wire \weights_inst.data_out[20] ;
 wire \weights_inst.data_out[21] ;
 wire \weights_inst.data_out[22] ;
 wire \weights_inst.data_out[23] ;
 wire \weights_inst.data_out[2] ;
 wire \weights_inst.data_out[3] ;
 wire \weights_inst.data_out[4] ;
 wire \weights_inst.data_out[5] ;
 wire \weights_inst.data_out[6] ;
 wire \weights_inst.data_out[7] ;
 wire \weights_inst.data_out[8] ;
 wire \weights_inst.data_out[9] ;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_0137_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(_0389_));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(_0424_));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(_0434_));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(_0449_));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(_0467_));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(_0560_));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(_0608_));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(_0617_));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(_0645_));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(_0645_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_0137_));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(_0725_));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(_0739_));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(_0764_));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(_0770_));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(_0787_));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(_0798_));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(_0840_));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(_0878_));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(_0888_));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(_0888_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_0177_));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(_0898_));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(_0900_));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(_0912_));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(_0926_));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(_0965_));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(_0965_));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(_0990_));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(_1001_));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(_1034_));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(_1038_));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_0204_));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(_1038_));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(_1038_));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(_1038_));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(_1038_));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(_1072_));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(_1088_));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(_1102_));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(_1103_));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(_1103_));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(_1154_));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_0215_));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(_1160_));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(_1173_));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(_1200_));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(_1200_));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(_1200_));
 sky130_fd_sc_hd__diode_2 ANTENNA_55 (.DIODE(_1202_));
 sky130_fd_sc_hd__diode_2 ANTENNA_56 (.DIODE(_1213_));
 sky130_fd_sc_hd__diode_2 ANTENNA_57 (.DIODE(_1253_));
 sky130_fd_sc_hd__diode_2 ANTENNA_58 (.DIODE(_1307_));
 sky130_fd_sc_hd__diode_2 ANTENNA_59 (.DIODE(_1354_));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_0253_));
 sky130_fd_sc_hd__diode_2 ANTENNA_60 (.DIODE(_1407_));
 sky130_fd_sc_hd__diode_2 ANTENNA_61 (.DIODE(_1407_));
 sky130_fd_sc_hd__diode_2 ANTENNA_62 (.DIODE(_1407_));
 sky130_fd_sc_hd__diode_2 ANTENNA_63 (.DIODE(_1407_));
 sky130_fd_sc_hd__diode_2 ANTENNA_64 (.DIODE(_1470_));
 sky130_fd_sc_hd__diode_2 ANTENNA_65 (.DIODE(_1482_));
 sky130_fd_sc_hd__diode_2 ANTENNA_66 (.DIODE(_1491_));
 sky130_fd_sc_hd__diode_2 ANTENNA_67 (.DIODE(_1494_));
 sky130_fd_sc_hd__diode_2 ANTENNA_68 (.DIODE(_0193_));
 sky130_fd_sc_hd__diode_2 ANTENNA_69 (.DIODE(_0733_));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(_0298_));
 sky130_fd_sc_hd__diode_2 ANTENNA_70 (.DIODE(_0764_));
 sky130_fd_sc_hd__diode_2 ANTENNA_71 (.DIODE(_0782_));
 sky130_fd_sc_hd__diode_2 ANTENNA_72 (.DIODE(_0782_));
 sky130_fd_sc_hd__diode_2 ANTENNA_73 (.DIODE(_0798_));
 sky130_fd_sc_hd__diode_2 ANTENNA_74 (.DIODE(_0798_));
 sky130_fd_sc_hd__diode_2 ANTENNA_75 (.DIODE(_0898_));
 sky130_fd_sc_hd__diode_2 ANTENNA_76 (.DIODE(_0900_));
 sky130_fd_sc_hd__diode_2 ANTENNA_77 (.DIODE(_0926_));
 sky130_fd_sc_hd__diode_2 ANTENNA_78 (.DIODE(_0948_));
 sky130_fd_sc_hd__diode_2 ANTENNA_79 (.DIODE(_1041_));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(_0340_));
 sky130_fd_sc_hd__diode_2 ANTENNA_80 (.DIODE(_1056_));
 sky130_fd_sc_hd__diode_2 ANTENNA_81 (.DIODE(_1063_));
 sky130_fd_sc_hd__diode_2 ANTENNA_82 (.DIODE(_1064_));
 sky130_fd_sc_hd__diode_2 ANTENNA_83 (.DIODE(_1190_));
 sky130_fd_sc_hd__diode_2 ANTENNA_84 (.DIODE(_1190_));
 sky130_fd_sc_hd__diode_2 ANTENNA_85 (.DIODE(_1265_));
 sky130_fd_sc_hd__diode_2 ANTENNA_86 (.DIODE(_1399_));
 sky130_fd_sc_hd__diode_2 ANTENNA_87 (.DIODE(_1064_));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(_0374_));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_331 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_448 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_395 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_31 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_336 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_366 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_303 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_506 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_196 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_525 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_395 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_525 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_284 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_310 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_170 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_339 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_89 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__nand2_1 _1533_ (.A(net17),
    .B(net12),
    .Y(_0420_));
 sky130_fd_sc_hd__nor2_1 _1534_ (.A(net87),
    .B(_0420_),
    .Y(_0003_));
 sky130_fd_sc_hd__xor2_4 _1535_ (.A(net7),
    .B(net9),
    .X(_0441_));
 sky130_fd_sc_hd__xor2_4 _1536_ (.A(net7),
    .B(net5),
    .X(_0452_));
 sky130_fd_sc_hd__and2_1 _1537_ (.A(net7),
    .B(net5),
    .X(_0462_));
 sky130_fd_sc_hd__a31o_4 _1538_ (.A1(net6),
    .A2(net4),
    .A3(net58),
    .B1(_0462_),
    .X(_0473_));
 sky130_fd_sc_hd__nand2_1 _1539_ (.A(net6),
    .B(net8),
    .Y(_0484_));
 sky130_fd_sc_hd__or2_1 _1540_ (.A(net6),
    .B(net8),
    .X(_0495_));
 sky130_fd_sc_hd__and2_2 _1541_ (.A(_0484_),
    .B(_0495_),
    .X(_0505_));
 sky130_fd_sc_hd__and3_4 _1542_ (.A(_0441_),
    .B(_0473_),
    .C(_0505_),
    .X(_0516_));
 sky130_fd_sc_hd__nand2_1 _1543_ (.A(net8),
    .B(net10),
    .Y(_0527_));
 sky130_fd_sc_hd__or2_2 _1544_ (.A(net8),
    .B(net10),
    .X(_0537_));
 sky130_fd_sc_hd__nand2_2 _1545_ (.A(_0527_),
    .B(_0537_),
    .Y(_0548_));
 sky130_fd_sc_hd__and2_1 _1546_ (.A(net7),
    .B(net9),
    .X(_0559_));
 sky130_fd_sc_hd__a31o_2 _1547_ (.A1(net6),
    .A2(net8),
    .A3(_0441_),
    .B1(_0559_),
    .X(_0570_));
 sky130_fd_sc_hd__xnor2_4 _1548_ (.A(_0548_),
    .B(_0570_),
    .Y(_0580_));
 sky130_fd_sc_hd__and2_1 _1549_ (.A(_0516_),
    .B(_0580_),
    .X(_0591_));
 sky130_fd_sc_hd__clkbuf_4 _1550_ (.A(_0591_),
    .X(_0602_));
 sky130_fd_sc_hd__a21boi_4 _1551_ (.A1(_0537_),
    .A2(_0570_),
    .B1_N(_0527_),
    .Y(_0613_));
 sky130_fd_sc_hd__xnor2_4 _1552_ (.A(net9),
    .B(_0613_),
    .Y(_0623_));
 sky130_fd_sc_hd__xnor2_4 _1553_ (.A(_0602_),
    .B(_0623_),
    .Y(_0634_));
 sky130_fd_sc_hd__buf_6 _1554_ (.A(_0634_),
    .X(_0645_));
 sky130_fd_sc_hd__clkbuf_4 _1555_ (.A(_0645_),
    .X(_0655_));
 sky130_fd_sc_hd__xor2_4 _1556_ (.A(_0516_),
    .B(_0580_),
    .X(_0661_));
 sky130_fd_sc_hd__clkbuf_8 _1557_ (.A(_0661_),
    .X(_0667_));
 sky130_fd_sc_hd__buf_4 _1558_ (.A(_0667_),
    .X(_0673_));
 sky130_fd_sc_hd__a21boi_4 _1559_ (.A1(_0473_),
    .A2(_0495_),
    .B1_N(_0484_),
    .Y(_0679_));
 sky130_fd_sc_hd__xor2_4 _1560_ (.A(_0441_),
    .B(_0679_),
    .X(_0685_));
 sky130_fd_sc_hd__buf_4 _1561_ (.A(_0685_),
    .X(_0694_));
 sky130_fd_sc_hd__buf_4 _1562_ (.A(_0694_),
    .X(_0703_));
 sky130_fd_sc_hd__buf_4 _1563_ (.A(_0703_),
    .X(_0706_));
 sky130_fd_sc_hd__buf_8 _1564_ (.A(net3),
    .X(_0708_));
 sky130_fd_sc_hd__xor2_4 _1565_ (.A(net6),
    .B(net4),
    .X(_0710_));
 sky130_fd_sc_hd__buf_12 _1566_ (.A(_0710_),
    .X(_0711_));
 sky130_fd_sc_hd__nand2_4 _1567_ (.A(_0708_),
    .B(_0711_),
    .Y(_0712_));
 sky130_fd_sc_hd__buf_4 _1568_ (.A(_0712_),
    .X(_0713_));
 sky130_fd_sc_hd__nand2_2 _1569_ (.A(net6),
    .B(net4),
    .Y(_0714_));
 sky130_fd_sc_hd__xor2_4 _1570_ (.A(net58),
    .B(_0714_),
    .X(_0715_));
 sky130_fd_sc_hd__buf_4 _1571_ (.A(_0715_),
    .X(_0716_));
 sky130_fd_sc_hd__clkbuf_8 _1572_ (.A(net2),
    .X(_0717_));
 sky130_fd_sc_hd__clkbuf_8 _1573_ (.A(_0717_),
    .X(_0718_));
 sky130_fd_sc_hd__nand2b_4 _1574_ (.A_N(net3),
    .B(_0718_),
    .Y(_0719_));
 sky130_fd_sc_hd__nor2_4 _1575_ (.A(_0711_),
    .B(_0719_),
    .Y(_0720_));
 sky130_fd_sc_hd__nor2_4 _1576_ (.A(_0716_),
    .B(_0720_),
    .Y(_0721_));
 sky130_fd_sc_hd__nand2_4 _1577_ (.A(_0713_),
    .B(_0721_),
    .Y(_0722_));
 sky130_fd_sc_hd__xnor2_4 _1578_ (.A(_0473_),
    .B(_0505_),
    .Y(_0723_));
 sky130_fd_sc_hd__buf_4 _1579_ (.A(_0723_),
    .X(_0724_));
 sky130_fd_sc_hd__buf_4 _1580_ (.A(_0724_),
    .X(_0725_));
 sky130_fd_sc_hd__xnor2_2 _1581_ (.A(net58),
    .B(_0714_),
    .Y(_0726_));
 sky130_fd_sc_hd__clkbuf_8 _1582_ (.A(_0726_),
    .X(_0727_));
 sky130_fd_sc_hd__buf_8 _1583_ (.A(_0727_),
    .X(_0728_));
 sky130_fd_sc_hd__inv_6 _1584_ (.A(net3),
    .Y(_0729_));
 sky130_fd_sc_hd__xnor2_4 _1585_ (.A(net6),
    .B(net4),
    .Y(_0730_));
 sky130_fd_sc_hd__buf_8 _1586_ (.A(_0730_),
    .X(_0731_));
 sky130_fd_sc_hd__nand2_4 _1587_ (.A(_0729_),
    .B(_0731_),
    .Y(_0732_));
 sky130_fd_sc_hd__nor2_8 _1588_ (.A(_0728_),
    .B(_0732_),
    .Y(_0733_));
 sky130_fd_sc_hd__nor2_2 _1589_ (.A(_0725_),
    .B(_0733_),
    .Y(_0734_));
 sky130_fd_sc_hd__clkbuf_16 _1590_ (.A(_0711_),
    .X(_0735_));
 sky130_fd_sc_hd__and2b_1 _1591_ (.A_N(net2),
    .B(net3),
    .X(_0736_));
 sky130_fd_sc_hd__buf_8 _1592_ (.A(_0736_),
    .X(_0737_));
 sky130_fd_sc_hd__nand2_4 _1593_ (.A(_0735_),
    .B(_0737_),
    .Y(_0738_));
 sky130_fd_sc_hd__clkbuf_8 _1594_ (.A(_0738_),
    .X(_0739_));
 sky130_fd_sc_hd__clkbuf_8 _1595_ (.A(_0727_),
    .X(_0740_));
 sky130_fd_sc_hd__clkbuf_8 _1596_ (.A(_0708_),
    .X(_0741_));
 sky130_fd_sc_hd__buf_8 _1597_ (.A(_0711_),
    .X(_0742_));
 sky130_fd_sc_hd__nor2_4 _1598_ (.A(_0741_),
    .B(_0742_),
    .Y(_0743_));
 sky130_fd_sc_hd__nor2_8 _1599_ (.A(_0740_),
    .B(_0743_),
    .Y(_0744_));
 sky130_fd_sc_hd__buf_4 _1600_ (.A(_0727_),
    .X(_0745_));
 sky130_fd_sc_hd__nand2_2 _1601_ (.A(_0718_),
    .B(_0731_),
    .Y(_0746_));
 sky130_fd_sc_hd__and3_2 _1602_ (.A(_0741_),
    .B(_0745_),
    .C(_0746_),
    .X(_0747_));
 sky130_fd_sc_hd__a21o_1 _1603_ (.A1(_0739_),
    .A2(_0744_),
    .B1(_0747_),
    .X(_0748_));
 sky130_fd_sc_hd__clkbuf_4 _1604_ (.A(_0723_),
    .X(_0749_));
 sky130_fd_sc_hd__buf_4 _1605_ (.A(_0749_),
    .X(_0750_));
 sky130_fd_sc_hd__buf_4 _1606_ (.A(_0750_),
    .X(_0751_));
 sky130_fd_sc_hd__clkbuf_4 _1607_ (.A(_0751_),
    .X(_0752_));
 sky130_fd_sc_hd__a22o_1 _1608_ (.A1(_0722_),
    .A2(_0734_),
    .B1(_0748_),
    .B2(_0752_),
    .X(_0753_));
 sky130_fd_sc_hd__clkbuf_8 _1609_ (.A(_0723_),
    .X(_0754_));
 sky130_fd_sc_hd__buf_6 _1610_ (.A(_0754_),
    .X(_0755_));
 sky130_fd_sc_hd__xnor2_4 _1611_ (.A(_0711_),
    .B(_0737_),
    .Y(_0756_));
 sky130_fd_sc_hd__clkbuf_8 _1612_ (.A(_0715_),
    .X(_0757_));
 sky130_fd_sc_hd__clkbuf_8 _1613_ (.A(_0757_),
    .X(_0758_));
 sky130_fd_sc_hd__and2b_1 _1614_ (.A_N(net3),
    .B(_0717_),
    .X(_0759_));
 sky130_fd_sc_hd__buf_8 _1615_ (.A(_0759_),
    .X(_0760_));
 sky130_fd_sc_hd__or3_4 _1616_ (.A(_0756_),
    .B(_0758_),
    .C(_0760_),
    .X(_0761_));
 sky130_fd_sc_hd__nand2_1 _1617_ (.A(_0755_),
    .B(_0761_),
    .Y(_0762_));
 sky130_fd_sc_hd__clkbuf_4 _1618_ (.A(_0715_),
    .X(_0763_));
 sky130_fd_sc_hd__and3_4 _1619_ (.A(_0763_),
    .B(_0719_),
    .C(_0712_),
    .X(_0764_));
 sky130_fd_sc_hd__clkbuf_16 _1620_ (.A(_0731_),
    .X(_0765_));
 sky130_fd_sc_hd__xnor2_4 _1621_ (.A(_0717_),
    .B(_0708_),
    .Y(_0766_));
 sky130_fd_sc_hd__nor2_8 _1622_ (.A(_0765_),
    .B(net57),
    .Y(_0767_));
 sky130_fd_sc_hd__buf_4 _1623_ (.A(_0715_),
    .X(_0768_));
 sky130_fd_sc_hd__clkbuf_8 _1624_ (.A(_0768_),
    .X(_0769_));
 sky130_fd_sc_hd__buf_6 _1625_ (.A(_0769_),
    .X(_0770_));
 sky130_fd_sc_hd__clkbuf_8 _1626_ (.A(_0765_),
    .X(_0771_));
 sky130_fd_sc_hd__buf_6 _1627_ (.A(_0718_),
    .X(_0772_));
 sky130_fd_sc_hd__a21oi_1 _1628_ (.A1(_0729_),
    .A2(_0771_),
    .B1(_0772_),
    .Y(_0773_));
 sky130_fd_sc_hd__nor2_2 _1629_ (.A(_0770_),
    .B(net52),
    .Y(_0774_));
 sky130_fd_sc_hd__nor2_2 _1630_ (.A(_0767_),
    .B(_0774_),
    .Y(_0775_));
 sky130_fd_sc_hd__xnor2_2 _1631_ (.A(_0441_),
    .B(_0679_),
    .Y(_0776_));
 sky130_fd_sc_hd__clkbuf_4 _1632_ (.A(_0776_),
    .X(_0777_));
 sky130_fd_sc_hd__clkbuf_8 _1633_ (.A(_0777_),
    .X(_0778_));
 sky130_fd_sc_hd__clkbuf_4 _1634_ (.A(_0778_),
    .X(_0779_));
 sky130_fd_sc_hd__o221a_1 _1635_ (.A1(_0762_),
    .A2(_0764_),
    .B1(_0775_),
    .B2(_0752_),
    .C1(_0779_),
    .X(_0780_));
 sky130_fd_sc_hd__a21oi_1 _1636_ (.A1(_0706_),
    .A2(_0753_),
    .B1(_0780_),
    .Y(_0781_));
 sky130_fd_sc_hd__clkbuf_8 _1637_ (.A(_0777_),
    .X(_0782_));
 sky130_fd_sc_hd__buf_4 _1638_ (.A(_0782_),
    .X(_0783_));
 sky130_fd_sc_hd__buf_8 _1639_ (.A(_0726_),
    .X(_0784_));
 sky130_fd_sc_hd__clkbuf_8 _1640_ (.A(_0784_),
    .X(_0785_));
 sky130_fd_sc_hd__buf_4 _1641_ (.A(_0785_),
    .X(_0786_));
 sky130_fd_sc_hd__nor2_8 _1642_ (.A(_0729_),
    .B(_0735_),
    .Y(_0787_));
 sky130_fd_sc_hd__nor2_8 _1643_ (.A(_0772_),
    .B(_0787_),
    .Y(_0788_));
 sky130_fd_sc_hd__o21a_1 _1644_ (.A1(_0786_),
    .A2(_0788_),
    .B1(_0755_),
    .X(_0789_));
 sky130_fd_sc_hd__nand2_4 _1645_ (.A(_0708_),
    .B(_0731_),
    .Y(_0790_));
 sky130_fd_sc_hd__nand2_4 _1646_ (.A(_0727_),
    .B(_0790_),
    .Y(_0791_));
 sky130_fd_sc_hd__nand2_1 _1647_ (.A(_0789_),
    .B(_0791_),
    .Y(_0792_));
 sky130_fd_sc_hd__or2b_1 _1648_ (.A(_0717_),
    .B_N(_0708_),
    .X(_0793_));
 sky130_fd_sc_hd__nand2_1 _1649_ (.A(_0742_),
    .B(_0793_),
    .Y(_0794_));
 sky130_fd_sc_hd__inv_2 _1650_ (.A(net2),
    .Y(_0795_));
 sky130_fd_sc_hd__nand2_2 _1651_ (.A(_0795_),
    .B(_0731_),
    .Y(_0796_));
 sky130_fd_sc_hd__buf_4 _1652_ (.A(_0796_),
    .X(_0797_));
 sky130_fd_sc_hd__and3_4 _1653_ (.A(_0794_),
    .B(_0728_),
    .C(_0797_),
    .X(_0798_));
 sky130_fd_sc_hd__buf_4 _1654_ (.A(_0723_),
    .X(_0799_));
 sky130_fd_sc_hd__clkbuf_8 _1655_ (.A(_0799_),
    .X(_0800_));
 sky130_fd_sc_hd__clkbuf_8 _1656_ (.A(_0800_),
    .X(_0801_));
 sky130_fd_sc_hd__buf_4 _1657_ (.A(_0732_),
    .X(_0802_));
 sky130_fd_sc_hd__buf_8 _1658_ (.A(_0802_),
    .X(_0803_));
 sky130_fd_sc_hd__nor2_1 _1659_ (.A(_0718_),
    .B(_0711_),
    .Y(_0804_));
 sky130_fd_sc_hd__clkbuf_8 _1660_ (.A(_0804_),
    .X(_0805_));
 sky130_fd_sc_hd__nor2_8 _1661_ (.A(_0740_),
    .B(_0805_),
    .Y(_0806_));
 sky130_fd_sc_hd__buf_4 _1662_ (.A(_0806_),
    .X(_0807_));
 sky130_fd_sc_hd__nand2_1 _1663_ (.A(_0803_),
    .B(_0807_),
    .Y(_0808_));
 sky130_fd_sc_hd__or3b_1 _1664_ (.A(_0798_),
    .B(_0801_),
    .C_N(_0808_),
    .X(_0809_));
 sky130_fd_sc_hd__buf_4 _1665_ (.A(_0799_),
    .X(_0810_));
 sky130_fd_sc_hd__buf_4 _1666_ (.A(_0810_),
    .X(_0811_));
 sky130_fd_sc_hd__nor2_1 _1667_ (.A(_0718_),
    .B(_0731_),
    .Y(_0812_));
 sky130_fd_sc_hd__clkbuf_8 _1668_ (.A(_0812_),
    .X(_0813_));
 sky130_fd_sc_hd__nor2_1 _1669_ (.A(_0768_),
    .B(_0813_),
    .Y(_0814_));
 sky130_fd_sc_hd__buf_4 _1670_ (.A(_0814_),
    .X(_0815_));
 sky130_fd_sc_hd__buf_4 _1671_ (.A(_0815_),
    .X(_0816_));
 sky130_fd_sc_hd__nand2_8 _1672_ (.A(_0765_),
    .B(_0766_),
    .Y(_0817_));
 sky130_fd_sc_hd__xnor2_2 _1673_ (.A(_0717_),
    .B(_0710_),
    .Y(_0818_));
 sky130_fd_sc_hd__clkbuf_8 _1674_ (.A(_0818_),
    .X(_0819_));
 sky130_fd_sc_hd__buf_4 _1675_ (.A(_0740_),
    .X(_0820_));
 sky130_fd_sc_hd__a21oi_1 _1676_ (.A1(_0713_),
    .A2(_0819_),
    .B1(_0820_),
    .Y(_0821_));
 sky130_fd_sc_hd__a21oi_1 _1677_ (.A1(_0816_),
    .A2(_0817_),
    .B1(_0821_),
    .Y(_0822_));
 sky130_fd_sc_hd__buf_4 _1678_ (.A(_0719_),
    .X(_0823_));
 sky130_fd_sc_hd__buf_4 _1679_ (.A(_0823_),
    .X(_0824_));
 sky130_fd_sc_hd__buf_6 _1680_ (.A(_0793_),
    .X(_0825_));
 sky130_fd_sc_hd__buf_4 _1681_ (.A(_0763_),
    .X(_0826_));
 sky130_fd_sc_hd__and3_4 _1682_ (.A(_0825_),
    .B(_0826_),
    .C(_0746_),
    .X(_0827_));
 sky130_fd_sc_hd__buf_8 _1683_ (.A(_0795_),
    .X(_0828_));
 sky130_fd_sc_hd__nand2_8 _1684_ (.A(_0828_),
    .B(_0742_),
    .Y(_0829_));
 sky130_fd_sc_hd__nand2_1 _1685_ (.A(_0717_),
    .B(_0708_),
    .Y(_0830_));
 sky130_fd_sc_hd__buf_4 _1686_ (.A(_0830_),
    .X(_0831_));
 sky130_fd_sc_hd__and4_2 _1687_ (.A(_0745_),
    .B(_0732_),
    .C(_0829_),
    .D(_0831_),
    .X(_0832_));
 sky130_fd_sc_hd__xor2_2 _1688_ (.A(_0473_),
    .B(_0505_),
    .X(_0833_));
 sky130_fd_sc_hd__clkbuf_4 _1689_ (.A(_0833_),
    .X(_0834_));
 sky130_fd_sc_hd__clkbuf_4 _1690_ (.A(_0834_),
    .X(_0835_));
 sky130_fd_sc_hd__buf_4 _1691_ (.A(_0835_),
    .X(_0836_));
 sky130_fd_sc_hd__a211o_1 _1692_ (.A1(_0824_),
    .A2(_0827_),
    .B1(_0832_),
    .C1(_0836_),
    .X(_0837_));
 sky130_fd_sc_hd__buf_4 _1693_ (.A(_0685_),
    .X(_0838_));
 sky130_fd_sc_hd__buf_4 _1694_ (.A(_0838_),
    .X(_0839_));
 sky130_fd_sc_hd__o211a_4 _1695_ (.A1(_0811_),
    .A2(_0822_),
    .B1(_0837_),
    .C1(_0839_),
    .X(_0840_));
 sky130_fd_sc_hd__xnor2_4 _1696_ (.A(_0516_),
    .B(_0580_),
    .Y(_0841_));
 sky130_fd_sc_hd__buf_4 _1697_ (.A(_0841_),
    .X(_0842_));
 sky130_fd_sc_hd__buf_4 _1698_ (.A(_0842_),
    .X(_0843_));
 sky130_fd_sc_hd__a311o_1 _1699_ (.A1(_0783_),
    .A2(_0792_),
    .A3(_0809_),
    .B1(_0840_),
    .C1(_0843_),
    .X(_0844_));
 sky130_fd_sc_hd__nand2_1 _1700_ (.A(_0602_),
    .B(_0623_),
    .Y(_0845_));
 sky130_fd_sc_hd__a31o_1 _1701_ (.A1(net8),
    .A2(net9),
    .A3(_0570_),
    .B1(net10),
    .X(_0846_));
 sky130_fd_sc_hd__nand3b_1 _1702_ (.A_N(_0613_),
    .B(net10),
    .C(net9),
    .Y(_0847_));
 sky130_fd_sc_hd__nand3_4 _1703_ (.A(_0845_),
    .B(net78),
    .C(net69),
    .Y(_0848_));
 sky130_fd_sc_hd__buf_8 _1704_ (.A(_0848_),
    .X(_0849_));
 sky130_fd_sc_hd__o211a_1 _1705_ (.A1(_0673_),
    .A2(_0781_),
    .B1(_0844_),
    .C1(_0849_),
    .X(_0850_));
 sky130_fd_sc_hd__nand2_4 _1706_ (.A(_0729_),
    .B(_0735_),
    .Y(_0851_));
 sky130_fd_sc_hd__nand2_8 _1707_ (.A(_0731_),
    .B(_0737_),
    .Y(_0852_));
 sky130_fd_sc_hd__nand2_1 _1708_ (.A(_0731_),
    .B(_0759_),
    .Y(_0853_));
 sky130_fd_sc_hd__clkbuf_8 _1709_ (.A(_0853_),
    .X(_0854_));
 sky130_fd_sc_hd__and3_4 _1710_ (.A(_0852_),
    .B(_0740_),
    .C(_0854_),
    .X(_0855_));
 sky130_fd_sc_hd__nand2_2 _1711_ (.A(_0851_),
    .B(_0855_),
    .Y(_0856_));
 sky130_fd_sc_hd__a21oi_1 _1712_ (.A1(_0808_),
    .A2(_0856_),
    .B1(_0849_),
    .Y(_0857_));
 sky130_fd_sc_hd__o21ai_1 _1713_ (.A1(net8),
    .A2(net9),
    .B1(net65),
    .Y(_0858_));
 sky130_fd_sc_hd__clkbuf_4 _1714_ (.A(net66),
    .X(_0859_));
 sky130_fd_sc_hd__xor2_4 _1715_ (.A(_0602_),
    .B(_0623_),
    .X(_0860_));
 sky130_fd_sc_hd__clkbuf_4 _1716_ (.A(_0860_),
    .X(_0861_));
 sky130_fd_sc_hd__and3_1 _1717_ (.A(_0845_),
    .B(_0846_),
    .C(_0847_),
    .X(_0862_));
 sky130_fd_sc_hd__clkbuf_4 _1718_ (.A(net70),
    .X(_0863_));
 sky130_fd_sc_hd__buf_4 _1719_ (.A(_0833_),
    .X(_0864_));
 sky130_fd_sc_hd__a21o_1 _1720_ (.A1(_0825_),
    .A2(_0769_),
    .B1(_0864_),
    .X(_0865_));
 sky130_fd_sc_hd__xnor2_4 _1721_ (.A(_0729_),
    .B(_0711_),
    .Y(_0866_));
 sky130_fd_sc_hd__buf_4 _1722_ (.A(_0866_),
    .X(_0867_));
 sky130_fd_sc_hd__nor2_8 _1723_ (.A(_0708_),
    .B(_0765_),
    .Y(_0868_));
 sky130_fd_sc_hd__nand2_1 _1724_ (.A(_0852_),
    .B(_0768_),
    .Y(_0869_));
 sky130_fd_sc_hd__a21o_1 _1725_ (.A1(_0718_),
    .A2(_0742_),
    .B1(_0741_),
    .X(_0870_));
 sky130_fd_sc_hd__or3b_4 _1726_ (.A(_0768_),
    .B(_0805_),
    .C_N(_0870_),
    .X(_0871_));
 sky130_fd_sc_hd__o21a_1 _1727_ (.A1(_0868_),
    .A2(_0869_),
    .B1(_0871_),
    .X(_0872_));
 sky130_fd_sc_hd__buf_4 _1728_ (.A(_0754_),
    .X(_0873_));
 sky130_fd_sc_hd__o32a_1 _1729_ (.A1(_0760_),
    .A2(_0865_),
    .A3(_0867_),
    .B1(_0872_),
    .B2(_0873_),
    .X(_0874_));
 sky130_fd_sc_hd__buf_4 _1730_ (.A(_0754_),
    .X(_0875_));
 sky130_fd_sc_hd__nand2_1 _1731_ (.A(_0815_),
    .B(_0817_),
    .Y(_0876_));
 sky130_fd_sc_hd__buf_6 _1732_ (.A(_0757_),
    .X(_0877_));
 sky130_fd_sc_hd__buf_6 _1733_ (.A(_0877_),
    .X(_0878_));
 sky130_fd_sc_hd__nand2_1 _1734_ (.A(_0878_),
    .B(_0813_),
    .Y(_0879_));
 sky130_fd_sc_hd__xnor2_4 _1735_ (.A(_0828_),
    .B(_0711_),
    .Y(_0880_));
 sky130_fd_sc_hd__buf_8 _1736_ (.A(_0729_),
    .X(_0881_));
 sky130_fd_sc_hd__nand2_2 _1737_ (.A(_0881_),
    .B(_0716_),
    .Y(_0882_));
 sky130_fd_sc_hd__and4_1 _1738_ (.A(_0864_),
    .B(_0823_),
    .C(_0880_),
    .D(_0882_),
    .X(_0883_));
 sky130_fd_sc_hd__a31o_1 _1739_ (.A1(_0875_),
    .A2(_0876_),
    .A3(_0879_),
    .B1(_0883_),
    .X(_0884_));
 sky130_fd_sc_hd__and2_1 _1740_ (.A(_0717_),
    .B(net3),
    .X(_0885_));
 sky130_fd_sc_hd__buf_6 _1741_ (.A(_0885_),
    .X(_0886_));
 sky130_fd_sc_hd__xnor2_4 _1742_ (.A(_0731_),
    .B(_0886_),
    .Y(_0887_));
 sky130_fd_sc_hd__nor2_4 _1743_ (.A(_0757_),
    .B(_0887_),
    .Y(_0888_));
 sky130_fd_sc_hd__or2_2 _1744_ (.A(_0864_),
    .B(_0888_),
    .X(_0889_));
 sky130_fd_sc_hd__nor2_8 _1745_ (.A(_0784_),
    .B(_0746_),
    .Y(_0890_));
 sky130_fd_sc_hd__or3_2 _1746_ (.A(_0717_),
    .B(_0708_),
    .C(_0710_),
    .X(_0891_));
 sky130_fd_sc_hd__buf_4 _1747_ (.A(_0891_),
    .X(_0892_));
 sky130_fd_sc_hd__nor2_2 _1748_ (.A(_0758_),
    .B(_0892_),
    .Y(_0893_));
 sky130_fd_sc_hd__a211o_1 _1749_ (.A1(_0806_),
    .A2(_0867_),
    .B1(_0893_),
    .C1(_0754_),
    .X(_0894_));
 sky130_fd_sc_hd__o21a_1 _1750_ (.A1(_0889_),
    .A2(_0890_),
    .B1(_0894_),
    .X(_0895_));
 sky130_fd_sc_hd__nor2_8 _1751_ (.A(_0717_),
    .B(_0708_),
    .Y(_0896_));
 sky130_fd_sc_hd__nand2_1 _1752_ (.A(_0742_),
    .B(_0896_),
    .Y(_0897_));
 sky130_fd_sc_hd__and3_2 _1753_ (.A(_0763_),
    .B(_0854_),
    .C(_0897_),
    .X(_0898_));
 sky130_fd_sc_hd__nor2_2 _1754_ (.A(_0772_),
    .B(_0768_),
    .Y(_0899_));
 sky130_fd_sc_hd__or2_4 _1755_ (.A(_0723_),
    .B(_0899_),
    .X(_0900_));
 sky130_fd_sc_hd__nor2_4 _1756_ (.A(_0828_),
    .B(_0765_),
    .Y(_0901_));
 sky130_fd_sc_hd__a32o_1 _1757_ (.A1(_0756_),
    .A2(_0768_),
    .A3(_0719_),
    .B1(_0813_),
    .B2(net58),
    .X(_0902_));
 sky130_fd_sc_hd__a21oi_4 _1758_ (.A1(_0741_),
    .A2(_0742_),
    .B1(_0718_),
    .Y(_0903_));
 sky130_fd_sc_hd__or2_1 _1759_ (.A(_0826_),
    .B(_0903_),
    .X(_0904_));
 sky130_fd_sc_hd__o221a_1 _1760_ (.A1(_0869_),
    .A2(_0901_),
    .B1(_0902_),
    .B2(_0799_),
    .C1(_0904_),
    .X(_0905_));
 sky130_fd_sc_hd__o21ba_1 _1761_ (.A1(_0898_),
    .A2(_0900_),
    .B1_N(_0905_),
    .X(_0906_));
 sky130_fd_sc_hd__buf_4 _1762_ (.A(_0661_),
    .X(_0907_));
 sky130_fd_sc_hd__mux4_1 _1763_ (.A0(_0874_),
    .A1(_0884_),
    .A2(_0895_),
    .A3(_0906_),
    .S0(_0782_),
    .S1(_0907_),
    .X(_0908_));
 sky130_fd_sc_hd__nor2_1 _1764_ (.A(_0863_),
    .B(_0908_),
    .Y(_0909_));
 sky130_fd_sc_hd__buf_4 _1765_ (.A(_0834_),
    .X(_0910_));
 sky130_fd_sc_hd__buf_4 _1766_ (.A(_0910_),
    .X(_0911_));
 sky130_fd_sc_hd__and3_2 _1767_ (.A(_0745_),
    .B(_0732_),
    .C(_0831_),
    .X(_0912_));
 sky130_fd_sc_hd__a21oi_4 _1768_ (.A1(_0881_),
    .A2(_0829_),
    .B1(_0785_),
    .Y(_0913_));
 sky130_fd_sc_hd__clkbuf_8 _1769_ (.A(_0776_),
    .X(_0914_));
 sky130_fd_sc_hd__buf_4 _1770_ (.A(_0914_),
    .X(_0915_));
 sky130_fd_sc_hd__buf_4 _1771_ (.A(_0790_),
    .X(_0916_));
 sky130_fd_sc_hd__buf_4 _1772_ (.A(_0916_),
    .X(_0917_));
 sky130_fd_sc_hd__clkbuf_8 _1773_ (.A(_0826_),
    .X(_0918_));
 sky130_fd_sc_hd__a21o_2 _1774_ (.A1(_0881_),
    .A2(_0819_),
    .B1(_0918_),
    .X(_0919_));
 sky130_fd_sc_hd__a21o_1 _1775_ (.A1(_0917_),
    .A2(_0919_),
    .B1(_0875_),
    .X(_0920_));
 sky130_fd_sc_hd__o311a_1 _1776_ (.A1(_0911_),
    .A2(_0912_),
    .A3(_0913_),
    .B1(_0915_),
    .C1(_0920_),
    .X(_0921_));
 sky130_fd_sc_hd__buf_6 _1777_ (.A(_0799_),
    .X(_0922_));
 sky130_fd_sc_hd__buf_4 _1778_ (.A(_0922_),
    .X(_0923_));
 sky130_fd_sc_hd__buf_4 _1779_ (.A(_0746_),
    .X(_0924_));
 sky130_fd_sc_hd__and3_4 _1780_ (.A(_0825_),
    .B(_0728_),
    .C(_0924_),
    .X(_0925_));
 sky130_fd_sc_hd__clkbuf_8 _1781_ (.A(_0757_),
    .X(_0926_));
 sky130_fd_sc_hd__nand2_1 _1782_ (.A(_0742_),
    .B(_0886_),
    .Y(_0927_));
 sky130_fd_sc_hd__and3_2 _1783_ (.A(_0926_),
    .B(_0802_),
    .C(_0927_),
    .X(_0928_));
 sky130_fd_sc_hd__buf_4 _1784_ (.A(_0851_),
    .X(_0929_));
 sky130_fd_sc_hd__nor2_4 _1785_ (.A(_0742_),
    .B(_0830_),
    .Y(_0930_));
 sky130_fd_sc_hd__nor2_8 _1786_ (.A(_0727_),
    .B(_0930_),
    .Y(_0931_));
 sky130_fd_sc_hd__a211o_1 _1787_ (.A1(_0788_),
    .A2(_0929_),
    .B1(_0931_),
    .C1(_0836_),
    .X(_0932_));
 sky130_fd_sc_hd__o311a_1 _1788_ (.A1(_0923_),
    .A2(_0925_),
    .A3(_0928_),
    .B1(_0932_),
    .C1(_0839_),
    .X(_0933_));
 sky130_fd_sc_hd__clkbuf_8 _1789_ (.A(_0777_),
    .X(_0934_));
 sky130_fd_sc_hd__buf_4 _1790_ (.A(_0934_),
    .X(_0935_));
 sky130_fd_sc_hd__buf_4 _1791_ (.A(_0910_),
    .X(_0936_));
 sky130_fd_sc_hd__nand2_4 _1792_ (.A(_0771_),
    .B(_0886_),
    .Y(_0937_));
 sky130_fd_sc_hd__and3_2 _1793_ (.A(_0918_),
    .B(_0738_),
    .C(_0937_),
    .X(_0938_));
 sky130_fd_sc_hd__clkbuf_4 _1794_ (.A(_0727_),
    .X(_0939_));
 sky130_fd_sc_hd__and3_4 _1795_ (.A(_0939_),
    .B(_0802_),
    .C(_0924_),
    .X(_0940_));
 sky130_fd_sc_hd__nor2_1 _1796_ (.A(_0758_),
    .B(_0866_),
    .Y(_0941_));
 sky130_fd_sc_hd__or2_2 _1797_ (.A(_0754_),
    .B(_0941_),
    .X(_0942_));
 sky130_fd_sc_hd__o32a_1 _1798_ (.A1(_0936_),
    .A2(_0938_),
    .A3(_0940_),
    .B1(net52),
    .B2(_0942_),
    .X(_0943_));
 sky130_fd_sc_hd__buf_4 _1799_ (.A(_0834_),
    .X(_0944_));
 sky130_fd_sc_hd__buf_4 _1800_ (.A(_0944_),
    .X(_0945_));
 sky130_fd_sc_hd__xnor2_4 _1801_ (.A(_0708_),
    .B(_0710_),
    .Y(_0946_));
 sky130_fd_sc_hd__buf_4 _1802_ (.A(_0897_),
    .X(_0947_));
 sky130_fd_sc_hd__nor2_8 _1803_ (.A(_0926_),
    .B(_0930_),
    .Y(_0948_));
 sky130_fd_sc_hd__nand2_1 _1804_ (.A(_0947_),
    .B(_0948_),
    .Y(_0949_));
 sky130_fd_sc_hd__buf_4 _1805_ (.A(_0685_),
    .X(_0950_));
 sky130_fd_sc_hd__a221o_1 _1806_ (.A1(_0945_),
    .A2(net56),
    .B1(_0882_),
    .B2(_0949_),
    .C1(_0950_),
    .X(_0951_));
 sky130_fd_sc_hd__buf_4 _1807_ (.A(_0842_),
    .X(_0952_));
 sky130_fd_sc_hd__o211ai_1 _1808_ (.A1(_0935_),
    .A2(_0943_),
    .B1(_0951_),
    .C1(_0952_),
    .Y(_0953_));
 sky130_fd_sc_hd__o311a_1 _1809_ (.A1(_0843_),
    .A2(_0921_),
    .A3(_0933_),
    .B1(_0953_),
    .C1(_0863_),
    .X(_0954_));
 sky130_fd_sc_hd__or3_1 _1810_ (.A(_0861_),
    .B(_0909_),
    .C(_0954_),
    .X(_0955_));
 sky130_fd_sc_hd__o311a_1 _1811_ (.A1(_0655_),
    .A2(_0850_),
    .A3(_0857_),
    .B1(_0859_),
    .C1(_0955_),
    .X(_0004_));
 sky130_fd_sc_hd__buf_4 _1812_ (.A(_0749_),
    .X(_0956_));
 sky130_fd_sc_hd__buf_4 _1813_ (.A(_0956_),
    .X(_0957_));
 sky130_fd_sc_hd__or2_1 _1814_ (.A(net2),
    .B(net3),
    .X(_0958_));
 sky130_fd_sc_hd__buf_4 _1815_ (.A(_0958_),
    .X(_0959_));
 sky130_fd_sc_hd__and3_2 _1816_ (.A(_0745_),
    .B(_0790_),
    .C(_0959_),
    .X(_0960_));
 sky130_fd_sc_hd__nand2_4 _1817_ (.A(_0771_),
    .B(_0959_),
    .Y(_0961_));
 sky130_fd_sc_hd__and2_1 _1818_ (.A(_0877_),
    .B(_0961_),
    .X(_0962_));
 sky130_fd_sc_hd__buf_4 _1819_ (.A(_0685_),
    .X(_0963_));
 sky130_fd_sc_hd__clkbuf_4 _1820_ (.A(_0834_),
    .X(_0964_));
 sky130_fd_sc_hd__a21o_4 _1821_ (.A1(_0729_),
    .A2(_0731_),
    .B1(_0795_),
    .X(_0965_));
 sky130_fd_sc_hd__and3_4 _1822_ (.A(_0716_),
    .B(_0796_),
    .C(_0965_),
    .X(_0966_));
 sky130_fd_sc_hd__and3_1 _1823_ (.A(_0784_),
    .B(_0719_),
    .C(_0790_),
    .X(_0967_));
 sky130_fd_sc_hd__or3_1 _1824_ (.A(_0964_),
    .B(_0966_),
    .C(_0967_),
    .X(_0968_));
 sky130_fd_sc_hd__o311a_1 _1825_ (.A1(_0957_),
    .A2(_0960_),
    .A3(_0962_),
    .B1(_0963_),
    .C1(_0968_),
    .X(_0969_));
 sky130_fd_sc_hd__buf_4 _1826_ (.A(_0926_),
    .X(_0970_));
 sky130_fd_sc_hd__buf_4 _1827_ (.A(_0797_),
    .X(_0971_));
 sky130_fd_sc_hd__nand2_1 _1828_ (.A(_0711_),
    .B(_0959_),
    .Y(_0972_));
 sky130_fd_sc_hd__clkbuf_8 _1829_ (.A(_0972_),
    .X(_0973_));
 sky130_fd_sc_hd__and3_2 _1830_ (.A(_0970_),
    .B(_0971_),
    .C(_0973_),
    .X(_0974_));
 sky130_fd_sc_hd__clkbuf_8 _1831_ (.A(_0939_),
    .X(_0975_));
 sky130_fd_sc_hd__nand2_8 _1832_ (.A(_0742_),
    .B(net57),
    .Y(_0976_));
 sky130_fd_sc_hd__and3_2 _1833_ (.A(_0975_),
    .B(_0971_),
    .C(_0976_),
    .X(_0977_));
 sky130_fd_sc_hd__buf_4 _1834_ (.A(_0777_),
    .X(_0978_));
 sky130_fd_sc_hd__nor2_1 _1835_ (.A(_0918_),
    .B(_0870_),
    .Y(_0979_));
 sky130_fd_sc_hd__nor2_2 _1836_ (.A(_0756_),
    .B(_0820_),
    .Y(_0980_));
 sky130_fd_sc_hd__or3_1 _1837_ (.A(_0944_),
    .B(_0979_),
    .C(_0980_),
    .X(_0981_));
 sky130_fd_sc_hd__o311a_1 _1838_ (.A1(_0751_),
    .A2(_0974_),
    .A3(_0977_),
    .B1(_0978_),
    .C1(_0981_),
    .X(_0982_));
 sky130_fd_sc_hd__buf_4 _1839_ (.A(_0959_),
    .X(_0983_));
 sky130_fd_sc_hd__buf_4 _1840_ (.A(_0833_),
    .X(_0984_));
 sky130_fd_sc_hd__clkbuf_8 _1841_ (.A(_0984_),
    .X(_0985_));
 sky130_fd_sc_hd__a221o_1 _1842_ (.A1(_0916_),
    .A2(_0815_),
    .B1(_0983_),
    .B2(_0931_),
    .C1(_0985_),
    .X(_0986_));
 sky130_fd_sc_hd__o21ai_1 _1843_ (.A1(_0898_),
    .A2(_0899_),
    .B1(_0936_),
    .Y(_0987_));
 sky130_fd_sc_hd__and3_4 _1844_ (.A(_0758_),
    .B(_0937_),
    .C(_0947_),
    .X(_0988_));
 sky130_fd_sc_hd__nand2_8 _1845_ (.A(_0742_),
    .B(_0831_),
    .Y(_0989_));
 sky130_fd_sc_hd__nor2_4 _1846_ (.A(_0740_),
    .B(_0896_),
    .Y(_0990_));
 sky130_fd_sc_hd__a311o_1 _1847_ (.A1(_0937_),
    .A2(_0989_),
    .A3(_0990_),
    .B1(_0967_),
    .C1(_0984_),
    .X(_0991_));
 sky130_fd_sc_hd__o311a_1 _1848_ (.A1(_0750_),
    .A2(_0925_),
    .A3(_0988_),
    .B1(_0991_),
    .C1(_0838_),
    .X(_0992_));
 sky130_fd_sc_hd__buf_4 _1849_ (.A(_0661_),
    .X(_0993_));
 sky130_fd_sc_hd__a311o_1 _1850_ (.A1(_0978_),
    .A2(_0986_),
    .A3(_0987_),
    .B1(_0992_),
    .C1(_0993_),
    .X(_0994_));
 sky130_fd_sc_hd__o311a_1 _1851_ (.A1(_0952_),
    .A2(_0969_),
    .A3(_0982_),
    .B1(_0994_),
    .C1(_0860_),
    .X(_0995_));
 sky130_fd_sc_hd__nand2_8 _1852_ (.A(_0718_),
    .B(_0711_),
    .Y(_0996_));
 sky130_fd_sc_hd__nor2_2 _1853_ (.A(_0758_),
    .B(_0996_),
    .Y(_0997_));
 sky130_fd_sc_hd__xor2_1 _1854_ (.A(_0717_),
    .B(net3),
    .X(_0998_));
 sky130_fd_sc_hd__buf_4 _1855_ (.A(_0998_),
    .X(_0999_));
 sky130_fd_sc_hd__buf_4 _1856_ (.A(_0999_),
    .X(_1000_));
 sky130_fd_sc_hd__nand2_4 _1857_ (.A(_0826_),
    .B(_0996_),
    .Y(_1001_));
 sky130_fd_sc_hd__nor2_1 _1858_ (.A(_1000_),
    .B(_1001_),
    .Y(_1002_));
 sky130_fd_sc_hd__clkbuf_8 _1859_ (.A(_0794_),
    .X(_1003_));
 sky130_fd_sc_hd__and2_1 _1860_ (.A(_1003_),
    .B(_0785_),
    .X(_1004_));
 sky130_fd_sc_hd__a211o_1 _1861_ (.A1(_0824_),
    .A2(_0807_),
    .B1(_1004_),
    .C1(_0836_),
    .X(_1005_));
 sky130_fd_sc_hd__o311a_1 _1862_ (.A1(_0923_),
    .A2(_0997_),
    .A3(_1002_),
    .B1(_0839_),
    .C1(_1005_),
    .X(_1006_));
 sky130_fd_sc_hd__nor2_4 _1863_ (.A(_0765_),
    .B(_0760_),
    .Y(_1007_));
 sky130_fd_sc_hd__a21o_1 _1864_ (.A1(_0820_),
    .A2(_1007_),
    .B1(_0984_),
    .X(_1008_));
 sky130_fd_sc_hd__and3_1 _1865_ (.A(_0877_),
    .B(_0738_),
    .C(_0817_),
    .X(_1009_));
 sky130_fd_sc_hd__or2_1 _1866_ (.A(_1008_),
    .B(_1009_),
    .X(_1010_));
 sky130_fd_sc_hd__buf_4 _1867_ (.A(_0785_),
    .X(_1011_));
 sky130_fd_sc_hd__nand2_2 _1868_ (.A(_0852_),
    .B(_1003_),
    .Y(_1012_));
 sky130_fd_sc_hd__clkbuf_8 _1869_ (.A(_0823_),
    .X(_1013_));
 sky130_fd_sc_hd__nand2_1 _1870_ (.A(_1012_),
    .B(_1013_),
    .Y(_1014_));
 sky130_fd_sc_hd__clkbuf_8 _1871_ (.A(_0784_),
    .X(_1015_));
 sky130_fd_sc_hd__nor2_4 _1872_ (.A(_0741_),
    .B(_1015_),
    .Y(_1016_));
 sky130_fd_sc_hd__a2111o_1 _1873_ (.A1(_1011_),
    .A2(_1014_),
    .B1(_1016_),
    .C1(_0890_),
    .D1(_0922_),
    .X(_1017_));
 sky130_fd_sc_hd__a31o_1 _1874_ (.A1(_0915_),
    .A2(_1010_),
    .A3(_1017_),
    .B1(_0993_),
    .X(_1018_));
 sky130_fd_sc_hd__buf_4 _1875_ (.A(_0713_),
    .X(_1019_));
 sky130_fd_sc_hd__buf_4 _1876_ (.A(_0831_),
    .X(_1020_));
 sky130_fd_sc_hd__a221o_1 _1877_ (.A1(_0786_),
    .A2(_1019_),
    .B1(_0807_),
    .B2(_1020_),
    .C1(_0755_),
    .X(_1021_));
 sky130_fd_sc_hd__nor2_2 _1878_ (.A(_1012_),
    .B(_0970_),
    .Y(_1022_));
 sky130_fd_sc_hd__nor2_4 _1879_ (.A(_0820_),
    .B(net52),
    .Y(_1023_));
 sky130_fd_sc_hd__o21ai_1 _1880_ (.A1(_1022_),
    .A2(_1023_),
    .B1(_0801_),
    .Y(_1024_));
 sky130_fd_sc_hd__nand2_4 _1881_ (.A(_0735_),
    .B(_0760_),
    .Y(_1025_));
 sky130_fd_sc_hd__and3_2 _1882_ (.A(_0740_),
    .B(_0796_),
    .C(_1025_),
    .X(_1026_));
 sky130_fd_sc_hd__and3_2 _1883_ (.A(_0763_),
    .B(_0796_),
    .C(_0946_),
    .X(_1027_));
 sky130_fd_sc_hd__clkbuf_8 _1884_ (.A(_0834_),
    .X(_1028_));
 sky130_fd_sc_hd__o21ai_1 _1885_ (.A1(_1026_),
    .A2(_1027_),
    .B1(_1028_),
    .Y(_1029_));
 sky130_fd_sc_hd__nor2_4 _1886_ (.A(_0745_),
    .B(_0760_),
    .Y(_1030_));
 sky130_fd_sc_hd__nor2_4 _1887_ (.A(_0795_),
    .B(_0710_),
    .Y(_1031_));
 sky130_fd_sc_hd__nor2_1 _1888_ (.A(_0763_),
    .B(_1031_),
    .Y(_1032_));
 sky130_fd_sc_hd__a211o_1 _1889_ (.A1(_0756_),
    .A2(_1030_),
    .B1(_1032_),
    .C1(_0864_),
    .X(_1033_));
 sky130_fd_sc_hd__a31o_1 _1890_ (.A1(_0694_),
    .A2(_1029_),
    .A3(_1033_),
    .B1(_0841_),
    .X(_1034_));
 sky130_fd_sc_hd__a31o_1 _1891_ (.A1(_0915_),
    .A2(_1021_),
    .A3(_1024_),
    .B1(_1034_),
    .X(_1035_));
 sky130_fd_sc_hd__buf_8 _1892_ (.A(_0634_),
    .X(_1036_));
 sky130_fd_sc_hd__o211a_1 _1893_ (.A1(_1006_),
    .A2(_1018_),
    .B1(_1035_),
    .C1(_1036_),
    .X(_1037_));
 sky130_fd_sc_hd__o21ai_4 _1894_ (.A1(_0995_),
    .A2(_1037_),
    .B1(_0849_),
    .Y(_1038_));
 sky130_fd_sc_hd__buf_4 _1895_ (.A(_0860_),
    .X(_1039_));
 sky130_fd_sc_hd__clkbuf_4 _1896_ (.A(_1028_),
    .X(_1040_));
 sky130_fd_sc_hd__buf_4 _1897_ (.A(_0826_),
    .X(_1041_));
 sky130_fd_sc_hd__and3_2 _1898_ (.A(_1041_),
    .B(_0996_),
    .C(_0892_),
    .X(_1042_));
 sky130_fd_sc_hd__buf_4 _1899_ (.A(_1032_),
    .X(_1043_));
 sky130_fd_sc_hd__nor2_4 _1900_ (.A(_0828_),
    .B(_0868_),
    .Y(_1044_));
 sky130_fd_sc_hd__nor2_2 _1901_ (.A(_1015_),
    .B(_1044_),
    .Y(_1045_));
 sky130_fd_sc_hd__a221o_1 _1902_ (.A1(_1019_),
    .A2(_1043_),
    .B1(_0916_),
    .B2(_1045_),
    .C1(_0800_),
    .X(_1046_));
 sky130_fd_sc_hd__clkbuf_8 _1903_ (.A(_0838_),
    .X(_1047_));
 sky130_fd_sc_hd__o311a_1 _1904_ (.A1(_1040_),
    .A2(_0774_),
    .A3(_1042_),
    .B1(_1046_),
    .C1(_1047_),
    .X(_1048_));
 sky130_fd_sc_hd__clkbuf_4 _1905_ (.A(_0864_),
    .X(_1049_));
 sky130_fd_sc_hd__nor2_4 _1906_ (.A(_1003_),
    .B(_1015_),
    .Y(_1050_));
 sky130_fd_sc_hd__or3_1 _1907_ (.A(_1049_),
    .B(_0979_),
    .C(_1050_),
    .X(_1051_));
 sky130_fd_sc_hd__nor2_2 _1908_ (.A(_0765_),
    .B(_0831_),
    .Y(_1052_));
 sky130_fd_sc_hd__nor2_2 _1909_ (.A(_0757_),
    .B(_1052_),
    .Y(_1053_));
 sky130_fd_sc_hd__nand2_2 _1910_ (.A(_0802_),
    .B(_1053_),
    .Y(_1054_));
 sky130_fd_sc_hd__nand2_4 _1911_ (.A(_0737_),
    .B(_0877_),
    .Y(_1055_));
 sky130_fd_sc_hd__clkbuf_8 _1912_ (.A(_0724_),
    .X(_1056_));
 sky130_fd_sc_hd__a21o_1 _1913_ (.A1(_1054_),
    .A2(_1055_),
    .B1(_1056_),
    .X(_1057_));
 sky130_fd_sc_hd__a21oi_1 _1914_ (.A1(_1051_),
    .A2(_1057_),
    .B1(_0703_),
    .Y(_1058_));
 sky130_fd_sc_hd__nor2_8 _1915_ (.A(_0728_),
    .B(_0901_),
    .Y(_1059_));
 sky130_fd_sc_hd__buf_4 _1916_ (.A(_0984_),
    .X(_1060_));
 sky130_fd_sc_hd__a211o_1 _1917_ (.A1(_0946_),
    .A2(_1059_),
    .B1(_1060_),
    .C1(_0832_),
    .X(_1061_));
 sky130_fd_sc_hd__a2111o_1 _1918_ (.A1(_1000_),
    .A2(_1043_),
    .B1(_1016_),
    .C1(_0890_),
    .D1(_0800_),
    .X(_1062_));
 sky130_fd_sc_hd__buf_8 _1919_ (.A(_0754_),
    .X(_1063_));
 sky130_fd_sc_hd__nor2_8 _1920_ (.A(_0735_),
    .B(_0999_),
    .Y(_1064_));
 sky130_fd_sc_hd__nand2_8 _1921_ (.A(_0926_),
    .B(_1064_),
    .Y(_1065_));
 sky130_fd_sc_hd__nor2_4 _1922_ (.A(_0784_),
    .B(_0767_),
    .Y(_1066_));
 sky130_fd_sc_hd__or3_4 _1923_ (.A(_0757_),
    .B(_0720_),
    .C(_1007_),
    .X(_1067_));
 sky130_fd_sc_hd__and3b_1 _1924_ (.A_N(_1066_),
    .B(_0864_),
    .C(_1067_),
    .X(_1068_));
 sky130_fd_sc_hd__a311oi_4 _1925_ (.A1(_1063_),
    .A2(_0722_),
    .A3(_1065_),
    .B1(_1068_),
    .C1(_0914_),
    .Y(_1069_));
 sky130_fd_sc_hd__a311o_1 _1926_ (.A1(_0782_),
    .A2(_1061_),
    .A3(_1062_),
    .B1(_1069_),
    .C1(_0993_),
    .X(_1070_));
 sky130_fd_sc_hd__o31a_1 _1927_ (.A1(_0952_),
    .A2(_1048_),
    .A3(_1058_),
    .B1(_1070_),
    .X(_1071_));
 sky130_fd_sc_hd__nor2_8 _1928_ (.A(_0784_),
    .B(_1031_),
    .Y(_1072_));
 sky130_fd_sc_hd__nand2_8 _1929_ (.A(_0765_),
    .B(net74),
    .Y(_1073_));
 sky130_fd_sc_hd__a221o_1 _1930_ (.A1(_0803_),
    .A2(_1072_),
    .B1(_1053_),
    .B2(_1073_),
    .C1(_1036_),
    .X(_1074_));
 sky130_fd_sc_hd__o211ai_1 _1931_ (.A1(_1039_),
    .A2(_1071_),
    .B1(net75),
    .C1(_0863_),
    .Y(_1075_));
 sky130_fd_sc_hd__and3_1 _1932_ (.A(net66),
    .B(_1038_),
    .C(_1075_),
    .X(_1076_));
 sky130_fd_sc_hd__clkbuf_1 _1933_ (.A(net76),
    .X(_0015_));
 sky130_fd_sc_hd__nor2_4 _1934_ (.A(_0757_),
    .B(_0901_),
    .Y(_1077_));
 sky130_fd_sc_hd__buf_6 _1935_ (.A(net57),
    .X(_1078_));
 sky130_fd_sc_hd__nor2_4 _1936_ (.A(_0939_),
    .B(_1078_),
    .Y(_1079_));
 sky130_fd_sc_hd__a221o_1 _1937_ (.A1(_0983_),
    .A2(_1077_),
    .B1(_1079_),
    .B2(_0971_),
    .C1(_0910_),
    .X(_1080_));
 sky130_fd_sc_hd__a211o_1 _1938_ (.A1(_0916_),
    .A2(_1045_),
    .B1(_0912_),
    .C1(_0724_),
    .X(_1081_));
 sky130_fd_sc_hd__nand2_1 _1939_ (.A(_1080_),
    .B(_1081_),
    .Y(_1082_));
 sky130_fd_sc_hd__buf_4 _1940_ (.A(_0799_),
    .X(_1083_));
 sky130_fd_sc_hd__nor2_4 _1941_ (.A(_0784_),
    .B(_0868_),
    .Y(_1084_));
 sky130_fd_sc_hd__nand2_1 _1942_ (.A(_0819_),
    .B(_1084_),
    .Y(_1085_));
 sky130_fd_sc_hd__a211oi_1 _1943_ (.A1(_0797_),
    .A2(_1084_),
    .B1(_0997_),
    .C1(_0754_),
    .Y(_1086_));
 sky130_fd_sc_hd__a31o_1 _1944_ (.A1(_1083_),
    .A2(_0856_),
    .A3(_1085_),
    .B1(_1086_),
    .X(_1087_));
 sky130_fd_sc_hd__nor2_4 _1945_ (.A(_0771_),
    .B(_0825_),
    .Y(_1088_));
 sky130_fd_sc_hd__buf_4 _1946_ (.A(_0772_),
    .X(_1089_));
 sky130_fd_sc_hd__nor2_1 _1947_ (.A(_0763_),
    .B(_0999_),
    .Y(_1090_));
 sky130_fd_sc_hd__or2_1 _1948_ (.A(_0723_),
    .B(_1090_),
    .X(_1091_));
 sky130_fd_sc_hd__a31o_1 _1949_ (.A1(_1089_),
    .A2(_0769_),
    .A3(_0713_),
    .B1(_1091_),
    .X(_1092_));
 sky130_fd_sc_hd__o41a_1 _1950_ (.A1(_0964_),
    .A2(_0760_),
    .A3(_1088_),
    .A4(_1059_),
    .B1(_1092_),
    .X(_1093_));
 sky130_fd_sc_hd__and3_2 _1951_ (.A(_0939_),
    .B(_0713_),
    .C(_0892_),
    .X(_1094_));
 sky130_fd_sc_hd__nand2_1 _1952_ (.A(_0802_),
    .B(_1072_),
    .Y(_1095_));
 sky130_fd_sc_hd__nand2_1 _1953_ (.A(_0724_),
    .B(_1095_),
    .Y(_1096_));
 sky130_fd_sc_hd__a21o_4 _1954_ (.A1(_0891_),
    .A2(_0973_),
    .B1(_0886_),
    .X(_1097_));
 sky130_fd_sc_hd__nand2_2 _1955_ (.A(_0769_),
    .B(_1097_),
    .Y(_1098_));
 sky130_fd_sc_hd__nor2_4 _1956_ (.A(_0757_),
    .B(_0767_),
    .Y(_1099_));
 sky130_fd_sc_hd__nor2_1 _1957_ (.A(_0754_),
    .B(_1099_),
    .Y(_1100_));
 sky130_fd_sc_hd__a2bb2o_1 _1958_ (.A1_N(_1094_),
    .A2_N(_1096_),
    .B1(_1098_),
    .B2(_1100_),
    .X(_1101_));
 sky130_fd_sc_hd__mux4_2 _1959_ (.A0(_1082_),
    .A1(_1087_),
    .A2(_1093_),
    .A3(_1101_),
    .S0(_0950_),
    .S1(_0842_),
    .X(_1102_));
 sky130_fd_sc_hd__and3_2 _1960_ (.A(_0852_),
    .B(_0785_),
    .C(_0823_),
    .X(_1103_));
 sky130_fd_sc_hd__nor2_1 _1961_ (.A(_1036_),
    .B(_1103_),
    .Y(_1104_));
 sky130_fd_sc_hd__nor2_1 _1962_ (.A(_0727_),
    .B(_0813_),
    .Y(_1105_));
 sky130_fd_sc_hd__buf_4 _1963_ (.A(_1105_),
    .X(_1106_));
 sky130_fd_sc_hd__nand2_2 _1964_ (.A(_0817_),
    .B(_1106_),
    .Y(_1107_));
 sky130_fd_sc_hd__a221o_1 _1965_ (.A1(_0645_),
    .A2(_1102_),
    .B1(_1104_),
    .B2(_1107_),
    .C1(_0848_),
    .X(_1108_));
 sky130_fd_sc_hd__buf_4 _1966_ (.A(_0944_),
    .X(_1109_));
 sky130_fd_sc_hd__nand2_2 _1967_ (.A(_0939_),
    .B(_0797_),
    .Y(_1110_));
 sky130_fd_sc_hd__nor2_2 _1968_ (.A(_0743_),
    .B(_1110_),
    .Y(_1111_));
 sky130_fd_sc_hd__and3_2 _1969_ (.A(_0826_),
    .B(_0829_),
    .C(_0831_),
    .X(_1112_));
 sky130_fd_sc_hd__nand2_2 _1970_ (.A(_0735_),
    .B(_0999_),
    .Y(_1113_));
 sky130_fd_sc_hd__a221o_1 _1971_ (.A1(_1113_),
    .A2(_1072_),
    .B1(_0929_),
    .B2(_0925_),
    .C1(_0750_),
    .X(_1114_));
 sky130_fd_sc_hd__buf_4 _1972_ (.A(_0838_),
    .X(_1115_));
 sky130_fd_sc_hd__o311a_1 _1973_ (.A1(_1109_),
    .A2(_1111_),
    .A3(_1112_),
    .B1(_1114_),
    .C1(_1115_),
    .X(_1116_));
 sky130_fd_sc_hd__buf_4 _1974_ (.A(_0745_),
    .X(_1117_));
 sky130_fd_sc_hd__nor2_1 _1975_ (.A(_1117_),
    .B(_0983_),
    .Y(_1118_));
 sky130_fd_sc_hd__nor2_1 _1976_ (.A(_0918_),
    .B(_0817_),
    .Y(_1119_));
 sky130_fd_sc_hd__nand2_2 _1977_ (.A(_0975_),
    .B(_1013_),
    .Y(_1120_));
 sky130_fd_sc_hd__a21o_1 _1978_ (.A1(_1120_),
    .A2(_0739_),
    .B1(_0836_),
    .X(_1121_));
 sky130_fd_sc_hd__o311a_1 _1979_ (.A1(_0751_),
    .A2(_1118_),
    .A3(_1119_),
    .B1(_0978_),
    .C1(_1121_),
    .X(_1122_));
 sky130_fd_sc_hd__clkbuf_8 _1980_ (.A(_0741_),
    .X(_1123_));
 sky130_fd_sc_hd__clkbuf_8 _1981_ (.A(_1123_),
    .X(_1124_));
 sky130_fd_sc_hd__nor2_2 _1982_ (.A(_0769_),
    .B(_0802_),
    .Y(_1125_));
 sky130_fd_sc_hd__a211o_1 _1983_ (.A1(_1124_),
    .A2(_1106_),
    .B1(_1125_),
    .C1(_1060_),
    .X(_1126_));
 sky130_fd_sc_hd__nor2_4 _1984_ (.A(_0826_),
    .B(net54),
    .Y(_1127_));
 sky130_fd_sc_hd__a311o_1 _1985_ (.A1(_0999_),
    .A2(_0916_),
    .A3(_1084_),
    .B1(_1127_),
    .C1(_0750_),
    .X(_1128_));
 sky130_fd_sc_hd__and3_2 _1986_ (.A(_0939_),
    .B(_0797_),
    .C(_0927_),
    .X(_1129_));
 sky130_fd_sc_hd__and3_2 _1987_ (.A(_0794_),
    .B(_0727_),
    .C(_0853_),
    .X(_1130_));
 sky130_fd_sc_hd__or3_1 _1988_ (.A(_0749_),
    .B(_1027_),
    .C(_1130_),
    .X(_1131_));
 sky130_fd_sc_hd__o311a_1 _1989_ (.A1(_0944_),
    .A2(_1066_),
    .A3(_1129_),
    .B1(_1131_),
    .C1(_0777_),
    .X(_1132_));
 sky130_fd_sc_hd__a311o_1 _1990_ (.A1(_1115_),
    .A2(_1126_),
    .A3(_1128_),
    .B1(_1132_),
    .C1(_0842_),
    .X(_1133_));
 sky130_fd_sc_hd__o311a_1 _1991_ (.A1(_0667_),
    .A2(_1116_),
    .A3(_1122_),
    .B1(_1133_),
    .C1(_0860_),
    .X(_1134_));
 sky130_fd_sc_hd__nor2_2 _1992_ (.A(_0881_),
    .B(_0786_),
    .Y(_1135_));
 sky130_fd_sc_hd__clkbuf_8 _1993_ (.A(_1015_),
    .X(_1136_));
 sky130_fd_sc_hd__and3_2 _1994_ (.A(_0716_),
    .B(_0738_),
    .C(_0796_),
    .X(_1137_));
 sky130_fd_sc_hd__a211o_1 _1995_ (.A1(_1136_),
    .A2(_0788_),
    .B1(_1137_),
    .C1(_1028_),
    .X(_1138_));
 sky130_fd_sc_hd__o21ai_1 _1996_ (.A1(_1091_),
    .A2(_1135_),
    .B1(_1138_),
    .Y(_1139_));
 sky130_fd_sc_hd__clkbuf_8 _1997_ (.A(_0984_),
    .X(_1140_));
 sky130_fd_sc_hd__nor2_2 _1998_ (.A(_0852_),
    .B(_1041_),
    .Y(_1141_));
 sky130_fd_sc_hd__nor2_1 _1999_ (.A(_1123_),
    .B(_1001_),
    .Y(_1142_));
 sky130_fd_sc_hd__and3_1 _2000_ (.A(_1003_),
    .B(_0926_),
    .C(_0823_),
    .X(_1143_));
 sky130_fd_sc_hd__o21ai_1 _2001_ (.A1(_0798_),
    .A2(_1143_),
    .B1(_1060_),
    .Y(_1144_));
 sky130_fd_sc_hd__o31a_1 _2002_ (.A1(_1140_),
    .A2(_1141_),
    .A3(_1142_),
    .B1(_1144_),
    .X(_1145_));
 sky130_fd_sc_hd__nand2_2 _2003_ (.A(_0828_),
    .B(_0758_),
    .Y(_1146_));
 sky130_fd_sc_hd__nand2_2 _2004_ (.A(_0835_),
    .B(_1146_),
    .Y(_1147_));
 sky130_fd_sc_hd__a21oi_1 _2005_ (.A1(_1013_),
    .A2(_1106_),
    .B1(_0925_),
    .Y(_1148_));
 sky130_fd_sc_hd__o32a_1 _2006_ (.A1(_1031_),
    .A2(_0868_),
    .A3(_1147_),
    .B1(_1148_),
    .B2(_0836_),
    .X(_1149_));
 sky130_fd_sc_hd__and3_2 _2007_ (.A(_0740_),
    .B(_0831_),
    .C(_0818_),
    .X(_1150_));
 sky130_fd_sc_hd__a31o_2 _2008_ (.A1(_0820_),
    .A2(_0823_),
    .A3(net54),
    .B1(_0799_),
    .X(_1151_));
 sky130_fd_sc_hd__and3_2 _2009_ (.A(_0716_),
    .B(_0924_),
    .C(_0851_),
    .X(_1152_));
 sky130_fd_sc_hd__o32a_1 _2010_ (.A1(_1140_),
    .A2(net52),
    .A3(_1150_),
    .B1(_1151_),
    .B2(_1152_),
    .X(_1153_));
 sky130_fd_sc_hd__mux4_2 _2011_ (.A0(_1139_),
    .A1(_1145_),
    .A2(_1149_),
    .A3(_1153_),
    .S0(_0778_),
    .S1(_0907_),
    .X(_1154_));
 sky130_fd_sc_hd__nor2_1 _2012_ (.A(_1039_),
    .B(_1154_),
    .Y(_1155_));
 sky130_fd_sc_hd__o21ai_1 _2013_ (.A1(_1134_),
    .A2(_1155_),
    .B1(_0849_),
    .Y(_1156_));
 sky130_fd_sc_hd__and3_1 _2014_ (.A(net66),
    .B(_1108_),
    .C(_1156_),
    .X(_1157_));
 sky130_fd_sc_hd__clkbuf_1 _2015_ (.A(net67),
    .X(_0019_));
 sky130_fd_sc_hd__clkbuf_4 _2016_ (.A(_0849_),
    .X(_1158_));
 sky130_fd_sc_hd__nor2_2 _2017_ (.A(_0741_),
    .B(_0812_),
    .Y(_1159_));
 sky130_fd_sc_hd__nand2_4 _2018_ (.A(_0975_),
    .B(_1159_),
    .Y(_1160_));
 sky130_fd_sc_hd__buf_4 _2019_ (.A(_1036_),
    .X(_1161_));
 sky130_fd_sc_hd__and3_2 _2020_ (.A(_0825_),
    .B(_0918_),
    .C(_0802_),
    .X(_1162_));
 sky130_fd_sc_hd__nor2_1 _2021_ (.A(_1161_),
    .B(_1162_),
    .Y(_1163_));
 sky130_fd_sc_hd__clkbuf_4 _2022_ (.A(_0993_),
    .X(_1164_));
 sky130_fd_sc_hd__buf_4 _2023_ (.A(_1049_),
    .X(_1165_));
 sky130_fd_sc_hd__nor2_2 _2024_ (.A(_1003_),
    .B(_0769_),
    .Y(_1166_));
 sky130_fd_sc_hd__nand2_4 _2025_ (.A(_0785_),
    .B(_0870_),
    .Y(_1167_));
 sky130_fd_sc_hd__nor2_2 _2026_ (.A(net58),
    .B(_0976_),
    .Y(_1168_));
 sky130_fd_sc_hd__nor2_1 _2027_ (.A(_0890_),
    .B(_1168_),
    .Y(_1169_));
 sky130_fd_sc_hd__a21o_1 _2028_ (.A1(_1167_),
    .A2(_1169_),
    .B1(_0725_),
    .X(_1170_));
 sky130_fd_sc_hd__o311a_1 _2029_ (.A1(_1165_),
    .A2(_1106_),
    .A3(_1166_),
    .B1(_1170_),
    .C1(_0703_),
    .X(_1171_));
 sky130_fd_sc_hd__nor2_2 _2030_ (.A(_0877_),
    .B(_1159_),
    .Y(_1172_));
 sky130_fd_sc_hd__a21o_4 _2031_ (.A1(_0772_),
    .A2(_0765_),
    .B1(_0741_),
    .X(_1173_));
 sky130_fd_sc_hd__nor2_2 _2032_ (.A(_1117_),
    .B(_1173_),
    .Y(_1174_));
 sky130_fd_sc_hd__nor2_4 _2033_ (.A(_0877_),
    .B(_1173_),
    .Y(_1175_));
 sky130_fd_sc_hd__nor2_1 _2034_ (.A(_0452_),
    .B(_0947_),
    .Y(_1176_));
 sky130_fd_sc_hd__or3_1 _2035_ (.A(_1049_),
    .B(_1175_),
    .C(_1176_),
    .X(_1177_));
 sky130_fd_sc_hd__buf_4 _2036_ (.A(_0914_),
    .X(_1178_));
 sky130_fd_sc_hd__o311a_1 _2037_ (.A1(_0811_),
    .A2(_1172_),
    .A3(_1174_),
    .B1(_1177_),
    .C1(_1178_),
    .X(_1179_));
 sky130_fd_sc_hd__buf_4 _2038_ (.A(_0750_),
    .X(_1180_));
 sky130_fd_sc_hd__nor2_4 _2039_ (.A(_0772_),
    .B(_0946_),
    .Y(_1181_));
 sky130_fd_sc_hd__nor2_2 _2040_ (.A(_0770_),
    .B(_1181_),
    .Y(_1182_));
 sky130_fd_sc_hd__nor2_4 _2041_ (.A(_0772_),
    .B(_1015_),
    .Y(_1183_));
 sky130_fd_sc_hd__and3_2 _2042_ (.A(_0745_),
    .B(_0887_),
    .C(_0959_),
    .X(_1184_));
 sky130_fd_sc_hd__or4_1 _2043_ (.A(_0835_),
    .B(_0733_),
    .C(_1183_),
    .D(_1184_),
    .X(_1185_));
 sky130_fd_sc_hd__o31ai_1 _2044_ (.A1(_1180_),
    .A2(_0756_),
    .A3(_1182_),
    .B1(_1185_),
    .Y(_1186_));
 sky130_fd_sc_hd__a31o_2 _2045_ (.A1(_0918_),
    .A2(_0823_),
    .A3(net54),
    .B1(_0864_),
    .X(_1187_));
 sky130_fd_sc_hd__nand2_2 _2046_ (.A(_0784_),
    .B(_0829_),
    .Y(_1188_));
 sky130_fd_sc_hd__nor2_2 _2047_ (.A(_1188_),
    .B(net56),
    .Y(_1189_));
 sky130_fd_sc_hd__nor2_8 _2048_ (.A(_0825_),
    .B(_0877_),
    .Y(_1190_));
 sky130_fd_sc_hd__nor2_1 _2049_ (.A(_0980_),
    .B(_1190_),
    .Y(_1191_));
 sky130_fd_sc_hd__o221a_1 _2050_ (.A1(_1187_),
    .A2(_1189_),
    .B1(_1191_),
    .B2(_0875_),
    .C1(_0914_),
    .X(_1192_));
 sky130_fd_sc_hd__buf_4 _2051_ (.A(_0841_),
    .X(_1193_));
 sky130_fd_sc_hd__a211o_1 _2052_ (.A1(_0703_),
    .A2(_1186_),
    .B1(_1192_),
    .C1(_1193_),
    .X(_1194_));
 sky130_fd_sc_hd__o31a_1 _2053_ (.A1(_1164_),
    .A2(_1171_),
    .A3(_1179_),
    .B1(_1194_),
    .X(_1195_));
 sky130_fd_sc_hd__o2bb2a_1 _2054_ (.A1_N(_1160_),
    .A2_N(_1163_),
    .B1(_1195_),
    .B2(_0861_),
    .X(_1196_));
 sky130_fd_sc_hd__clkbuf_4 _2055_ (.A(_0848_),
    .X(_1197_));
 sky130_fd_sc_hd__clkbuf_4 _2056_ (.A(_0934_),
    .X(_1198_));
 sky130_fd_sc_hd__buf_4 _2057_ (.A(_1041_),
    .X(_1199_));
 sky130_fd_sc_hd__and3_4 _2058_ (.A(_0852_),
    .B(_1015_),
    .C(_0851_),
    .X(_1200_));
 sky130_fd_sc_hd__a211o_1 _2059_ (.A1(_1199_),
    .A2(_1014_),
    .B1(_1200_),
    .C1(_1056_),
    .X(_1201_));
 sky130_fd_sc_hd__and2_4 _2060_ (.A(_0768_),
    .B(_0989_),
    .X(_1202_));
 sky130_fd_sc_hd__a211o_1 _2061_ (.A1(_1000_),
    .A2(_0816_),
    .B1(_1202_),
    .C1(_0945_),
    .X(_1203_));
 sky130_fd_sc_hd__nor2_2 _2062_ (.A(_0735_),
    .B(_0793_),
    .Y(_1204_));
 sky130_fd_sc_hd__nor2_1 _2063_ (.A(_1204_),
    .B(_0740_),
    .Y(_1205_));
 sky130_fd_sc_hd__clkbuf_8 _2064_ (.A(_1205_),
    .X(_1206_));
 sky130_fd_sc_hd__a211o_1 _2065_ (.A1(_0803_),
    .A2(_0815_),
    .B1(_1137_),
    .C1(_0964_),
    .X(_1207_));
 sky130_fd_sc_hd__o311a_1 _2066_ (.A1(_0875_),
    .A2(_1206_),
    .A3(_1094_),
    .B1(_1207_),
    .C1(_0950_),
    .X(_1208_));
 sky130_fd_sc_hd__a31o_1 _2067_ (.A1(_1198_),
    .A2(_1201_),
    .A3(_1203_),
    .B1(_1208_),
    .X(_1209_));
 sky130_fd_sc_hd__or4_1 _2068_ (.A(_0881_),
    .B(_0800_),
    .C(_0805_),
    .D(_1077_),
    .X(_1210_));
 sky130_fd_sc_hd__buf_4 _2069_ (.A(_0835_),
    .X(_1211_));
 sky130_fd_sc_hd__a221o_1 _2070_ (.A1(_0824_),
    .A2(_0815_),
    .B1(_1097_),
    .B2(_1199_),
    .C1(_1211_),
    .X(_1212_));
 sky130_fd_sc_hd__and2_4 _2071_ (.A(_0887_),
    .B(_0959_),
    .X(_1213_));
 sky130_fd_sc_hd__or3_2 _2072_ (.A(_0784_),
    .B(_0743_),
    .C(_0903_),
    .X(_1214_));
 sky130_fd_sc_hd__nor2_1 _2073_ (.A(net54),
    .B(_0868_),
    .Y(_1215_));
 sky130_fd_sc_hd__a221o_1 _2074_ (.A1(_1041_),
    .A2(_1213_),
    .B1(_1214_),
    .B2(_1215_),
    .C1(_0910_),
    .X(_1216_));
 sky130_fd_sc_hd__o311a_1 _2075_ (.A1(_1063_),
    .A2(_1099_),
    .A3(_1152_),
    .B1(_1216_),
    .C1(_0950_),
    .X(_1217_));
 sky130_fd_sc_hd__a31o_1 _2076_ (.A1(_1178_),
    .A2(_1210_),
    .A3(_1212_),
    .B1(_1217_),
    .X(_1218_));
 sky130_fd_sc_hd__buf_4 _2077_ (.A(_0924_),
    .X(_1219_));
 sky130_fd_sc_hd__nor2_1 _2078_ (.A(_0944_),
    .B(_1016_),
    .Y(_1220_));
 sky130_fd_sc_hd__nor2_4 _2079_ (.A(_0757_),
    .B(_0804_),
    .Y(_1221_));
 sky130_fd_sc_hd__a21o_1 _2080_ (.A1(_0739_),
    .A2(_1221_),
    .B1(_1168_),
    .X(_1222_));
 sky130_fd_sc_hd__a32o_1 _2081_ (.A1(_1019_),
    .A2(_1219_),
    .A3(_1220_),
    .B1(_1222_),
    .B2(_1211_),
    .X(_1223_));
 sky130_fd_sc_hd__and3_1 _2082_ (.A(_0828_),
    .B(_0763_),
    .C(_0866_),
    .X(_1224_));
 sky130_fd_sc_hd__or2_2 _2083_ (.A(_0834_),
    .B(_1224_),
    .X(_1225_));
 sky130_fd_sc_hd__or3b_1 _2084_ (.A(_1184_),
    .B(_0724_),
    .C_N(_1055_),
    .X(_1226_));
 sky130_fd_sc_hd__o21ai_1 _2085_ (.A1(_1044_),
    .A2(_1225_),
    .B1(_1226_),
    .Y(_1227_));
 sky130_fd_sc_hd__mux2_1 _2086_ (.A0(_1223_),
    .A1(_1227_),
    .S(_0839_),
    .X(_1228_));
 sky130_fd_sc_hd__buf_4 _2087_ (.A(_1221_),
    .X(_1229_));
 sky130_fd_sc_hd__and3_2 _2088_ (.A(_0926_),
    .B(_0738_),
    .C(_0924_),
    .X(_1230_));
 sky130_fd_sc_hd__a211o_1 _2089_ (.A1(_1229_),
    .A2(_1020_),
    .B1(_1230_),
    .C1(_0945_),
    .X(_1231_));
 sky130_fd_sc_hd__buf_4 _2090_ (.A(_0825_),
    .X(_1232_));
 sky130_fd_sc_hd__and3_1 _2091_ (.A(_1232_),
    .B(_0918_),
    .C(_0851_),
    .X(_1233_));
 sky130_fd_sc_hd__or2_1 _2092_ (.A(_0942_),
    .B(_1233_),
    .X(_1234_));
 sky130_fd_sc_hd__clkbuf_4 _2093_ (.A(_0835_),
    .X(_1235_));
 sky130_fd_sc_hd__nor2_4 _2094_ (.A(_0828_),
    .B(_0866_),
    .Y(_1236_));
 sky130_fd_sc_hd__a211o_1 _2095_ (.A1(_0929_),
    .A2(_0960_),
    .B1(_1236_),
    .C1(_0956_),
    .X(_1237_));
 sky130_fd_sc_hd__o311a_1 _2096_ (.A1(_1235_),
    .A2(_0912_),
    .A3(_0980_),
    .B1(_1237_),
    .C1(_0950_),
    .X(_1238_));
 sky130_fd_sc_hd__a31o_1 _2097_ (.A1(_1198_),
    .A2(_1231_),
    .A3(_1234_),
    .B1(_1238_),
    .X(_1239_));
 sky130_fd_sc_hd__mux4_2 _2098_ (.A0(_1209_),
    .A1(_1218_),
    .A2(_1228_),
    .A3(_1239_),
    .S0(_0843_),
    .S1(_1161_),
    .X(_1240_));
 sky130_fd_sc_hd__nand2_1 _2099_ (.A(_1197_),
    .B(_1240_),
    .Y(_1241_));
 sky130_fd_sc_hd__buf_2 _2100_ (.A(net66),
    .X(_1242_));
 sky130_fd_sc_hd__o211a_1 _2101_ (.A1(_1158_),
    .A2(_1196_),
    .B1(_1241_),
    .C1(_1242_),
    .X(_0021_));
 sky130_fd_sc_hd__buf_4 _2102_ (.A(_1193_),
    .X(_1243_));
 sky130_fd_sc_hd__buf_4 _2103_ (.A(_1040_),
    .X(_1244_));
 sky130_fd_sc_hd__a21oi_1 _2104_ (.A1(_1123_),
    .A2(_0971_),
    .B1(_0970_),
    .Y(_1245_));
 sky130_fd_sc_hd__nor2_2 _2105_ (.A(_1233_),
    .B(_1245_),
    .Y(_1246_));
 sky130_fd_sc_hd__and2_4 _2106_ (.A(_0763_),
    .B(_0891_),
    .X(_1247_));
 sky130_fd_sc_hd__or2_1 _2107_ (.A(_0810_),
    .B(_1247_),
    .X(_1248_));
 sky130_fd_sc_hd__nor2_4 _2108_ (.A(_1204_),
    .B(_0758_),
    .Y(_1249_));
 sky130_fd_sc_hd__clkbuf_4 _2109_ (.A(_0915_),
    .X(_1250_));
 sky130_fd_sc_hd__o221a_1 _2110_ (.A1(_1244_),
    .A2(_1246_),
    .B1(_1248_),
    .B2(_1249_),
    .C1(_1250_),
    .X(_1251_));
 sky130_fd_sc_hd__nor2_2 _2111_ (.A(_0826_),
    .B(_1064_),
    .Y(_1252_));
 sky130_fd_sc_hd__or2_4 _2112_ (.A(_0799_),
    .B(_1252_),
    .X(_1253_));
 sky130_fd_sc_hd__nand2_1 _2113_ (.A(_1123_),
    .B(_0924_),
    .Y(_1254_));
 sky130_fd_sc_hd__nor2_1 _2114_ (.A(_1136_),
    .B(_1254_),
    .Y(_1255_));
 sky130_fd_sc_hd__buf_4 _2115_ (.A(_0836_),
    .X(_1256_));
 sky130_fd_sc_hd__a211o_1 _2116_ (.A1(_1124_),
    .A2(_0816_),
    .B1(_1255_),
    .C1(_1256_),
    .X(_1257_));
 sky130_fd_sc_hd__o211a_1 _2117_ (.A1(_1183_),
    .A2(_1253_),
    .B1(_1257_),
    .C1(_0706_),
    .X(_1258_));
 sky130_fd_sc_hd__o21ai_4 _2118_ (.A1(_0786_),
    .A2(_0788_),
    .B1(_1063_),
    .Y(_1259_));
 sky130_fd_sc_hd__a21o_1 _2119_ (.A1(_1019_),
    .A2(_1043_),
    .B1(_1259_),
    .X(_1260_));
 sky130_fd_sc_hd__buf_4 _2120_ (.A(_1083_),
    .X(_1261_));
 sky130_fd_sc_hd__nor2_1 _2121_ (.A(_1261_),
    .B(_0938_),
    .Y(_1262_));
 sky130_fd_sc_hd__o21ai_1 _2122_ (.A1(_0791_),
    .A2(_1044_),
    .B1(_1262_),
    .Y(_1263_));
 sky130_fd_sc_hd__buf_4 _2123_ (.A(_0985_),
    .X(_1264_));
 sky130_fd_sc_hd__and3_4 _2124_ (.A(_0718_),
    .B(_0727_),
    .C(_0946_),
    .X(_1265_));
 sky130_fd_sc_hd__a21oi_1 _2125_ (.A1(_1123_),
    .A2(_0819_),
    .B1(_0975_),
    .Y(_1266_));
 sky130_fd_sc_hd__nor2_1 _2126_ (.A(_1117_),
    .B(_0916_),
    .Y(_1267_));
 sky130_fd_sc_hd__a311o_1 _2127_ (.A1(_1011_),
    .A2(_0739_),
    .A3(_0937_),
    .B1(_1267_),
    .C1(_1083_),
    .X(_1268_));
 sky130_fd_sc_hd__o311a_1 _2128_ (.A1(_1264_),
    .A2(_1265_),
    .A3(_1266_),
    .B1(_1268_),
    .C1(_1047_),
    .X(_1269_));
 sky130_fd_sc_hd__a31o_1 _2129_ (.A1(_0783_),
    .A2(_1260_),
    .A3(_1263_),
    .B1(_1269_),
    .X(_1270_));
 sky130_fd_sc_hd__nand2_1 _2130_ (.A(_1243_),
    .B(_1270_),
    .Y(_1271_));
 sky130_fd_sc_hd__o311a_1 _2131_ (.A1(_1243_),
    .A2(_1251_),
    .A3(_1258_),
    .B1(_1271_),
    .C1(_0655_),
    .X(_1272_));
 sky130_fd_sc_hd__clkbuf_4 _2132_ (.A(_1193_),
    .X(_1273_));
 sky130_fd_sc_hd__buf_4 _2133_ (.A(_0875_),
    .X(_1274_));
 sky130_fd_sc_hd__nand2_4 _2134_ (.A(_0745_),
    .B(_0712_),
    .Y(_1275_));
 sky130_fd_sc_hd__nor2_2 _2135_ (.A(_0760_),
    .B(_1275_),
    .Y(_1276_));
 sky130_fd_sc_hd__and3_4 _2136_ (.A(_0716_),
    .B(_0866_),
    .C(_0959_),
    .X(_1277_));
 sky130_fd_sc_hd__buf_4 _2137_ (.A(_0950_),
    .X(_1278_));
 sky130_fd_sc_hd__a211o_1 _2138_ (.A1(_0828_),
    .A2(_1084_),
    .B1(_1184_),
    .C1(_1264_),
    .X(_1279_));
 sky130_fd_sc_hd__o311a_1 _2139_ (.A1(_1274_),
    .A2(_1276_),
    .A3(_1277_),
    .B1(_1278_),
    .C1(_1279_),
    .X(_1280_));
 sky130_fd_sc_hd__buf_4 _2140_ (.A(_1109_),
    .X(_1281_));
 sky130_fd_sc_hd__and3_1 _2141_ (.A(_1232_),
    .B(_0770_),
    .C(_0854_),
    .X(_1282_));
 sky130_fd_sc_hd__nor2_1 _2142_ (.A(_0805_),
    .B(_1275_),
    .Y(_1283_));
 sky130_fd_sc_hd__or3b_1 _2143_ (.A(_1283_),
    .B(_0725_),
    .C_N(_1055_),
    .X(_1284_));
 sky130_fd_sc_hd__buf_4 _2144_ (.A(_0978_),
    .X(_1285_));
 sky130_fd_sc_hd__o311a_1 _2145_ (.A1(_1281_),
    .A2(_1265_),
    .A3(_1282_),
    .B1(_1284_),
    .C1(_1285_),
    .X(_1286_));
 sky130_fd_sc_hd__clkbuf_4 _2146_ (.A(_0963_),
    .X(_1287_));
 sky130_fd_sc_hd__and3_2 _2147_ (.A(_1117_),
    .B(_0854_),
    .C(_0927_),
    .X(_1288_));
 sky130_fd_sc_hd__a21oi_1 _2148_ (.A1(_1123_),
    .A2(_0971_),
    .B1(_1136_),
    .Y(_1289_));
 sky130_fd_sc_hd__o32a_1 _2149_ (.A1(_0725_),
    .A2(_1288_),
    .A3(_1289_),
    .B1(_1022_),
    .B2(_1187_),
    .X(_1290_));
 sky130_fd_sc_hd__buf_4 _2150_ (.A(_1063_),
    .X(_1291_));
 sky130_fd_sc_hd__a21oi_2 _2151_ (.A1(_0881_),
    .A2(_0819_),
    .B1(_0820_),
    .Y(_1292_));
 sky130_fd_sc_hd__a21oi_1 _2152_ (.A1(_1291_),
    .A2(_1292_),
    .B1(_0703_),
    .Y(_1293_));
 sky130_fd_sc_hd__and2_4 _2153_ (.A(_1015_),
    .B(_0887_),
    .X(_1294_));
 sky130_fd_sc_hd__a211o_1 _2154_ (.A1(_0971_),
    .A2(_1079_),
    .B1(_1294_),
    .C1(_0751_),
    .X(_1295_));
 sky130_fd_sc_hd__a221o_1 _2155_ (.A1(_1287_),
    .A2(_1290_),
    .B1(_1293_),
    .B2(_1295_),
    .C1(_0667_),
    .X(_1296_));
 sky130_fd_sc_hd__o311a_1 _2156_ (.A1(_1273_),
    .A2(_1280_),
    .A3(_1286_),
    .B1(_1296_),
    .C1(_1161_),
    .X(_1297_));
 sky130_fd_sc_hd__buf_4 _2157_ (.A(_1193_),
    .X(_1298_));
 sky130_fd_sc_hd__nand2_4 _2158_ (.A(_0755_),
    .B(_0882_),
    .Y(_1299_));
 sky130_fd_sc_hd__nor2_2 _2159_ (.A(_0878_),
    .B(_0961_),
    .Y(_1300_));
 sky130_fd_sc_hd__nor2_2 _2160_ (.A(net58),
    .B(_0771_),
    .Y(_1301_));
 sky130_fd_sc_hd__and2_2 _2161_ (.A(_1089_),
    .B(_1301_),
    .X(_1302_));
 sky130_fd_sc_hd__a221o_1 _2162_ (.A1(_1000_),
    .A2(_1043_),
    .B1(_1020_),
    .B2(_1301_),
    .C1(_1180_),
    .X(_1303_));
 sky130_fd_sc_hd__o311a_1 _2163_ (.A1(_1299_),
    .A2(_1300_),
    .A3(_1302_),
    .B1(_1303_),
    .C1(_0779_),
    .X(_1304_));
 sky130_fd_sc_hd__nor2_2 _2164_ (.A(_0826_),
    .B(_0989_),
    .Y(_1305_));
 sky130_fd_sc_hd__a21oi_1 _2165_ (.A1(_0891_),
    .A2(_0972_),
    .B1(_0768_),
    .Y(_1306_));
 sky130_fd_sc_hd__or3b_4 _2166_ (.A(_1306_),
    .B(_1056_),
    .C_N(_1107_),
    .X(_1307_));
 sky130_fd_sc_hd__buf_4 _2167_ (.A(_1115_),
    .X(_1308_));
 sky130_fd_sc_hd__o311a_1 _2168_ (.A1(_1281_),
    .A2(_0988_),
    .A3(_1305_),
    .B1(_1307_),
    .C1(_1308_),
    .X(_1309_));
 sky130_fd_sc_hd__clkbuf_4 _2169_ (.A(_1115_),
    .X(_1310_));
 sky130_fd_sc_hd__buf_4 _2170_ (.A(_0970_),
    .X(_1311_));
 sky130_fd_sc_hd__a221o_1 _2171_ (.A1(_1311_),
    .A2(_1064_),
    .B1(_1190_),
    .B2(_0945_),
    .C1(_0977_),
    .X(_1312_));
 sky130_fd_sc_hd__or4_1 _2172_ (.A(_0755_),
    .B(_1232_),
    .C(_1199_),
    .D(_0805_),
    .X(_1313_));
 sky130_fd_sc_hd__nor2_4 _2173_ (.A(_0735_),
    .B(_0785_),
    .Y(_1314_));
 sky130_fd_sc_hd__a21oi_1 _2174_ (.A1(_1123_),
    .A2(_0819_),
    .B1(_1041_),
    .Y(_1315_));
 sky130_fd_sc_hd__a211o_1 _2175_ (.A1(_0824_),
    .A2(_1314_),
    .B1(_1315_),
    .C1(_0985_),
    .X(_1316_));
 sky130_fd_sc_hd__o311a_1 _2176_ (.A1(_0957_),
    .A2(_1103_),
    .A3(_1255_),
    .B1(_1316_),
    .C1(_0778_),
    .X(_1317_));
 sky130_fd_sc_hd__clkbuf_8 _2177_ (.A(_0993_),
    .X(_1318_));
 sky130_fd_sc_hd__a311o_1 _2178_ (.A1(_1310_),
    .A2(_1312_),
    .A3(_1313_),
    .B1(_1317_),
    .C1(_1318_),
    .X(_1319_));
 sky130_fd_sc_hd__o311a_1 _2179_ (.A1(_1298_),
    .A2(_1304_),
    .A3(_1309_),
    .B1(_1319_),
    .C1(_1039_),
    .X(_1320_));
 sky130_fd_sc_hd__o21ai_1 _2180_ (.A1(_1297_),
    .A2(_1320_),
    .B1(_1197_),
    .Y(_1321_));
 sky130_fd_sc_hd__o311a_1 _2181_ (.A1(_1158_),
    .A2(_1163_),
    .A3(_1272_),
    .B1(_1321_),
    .C1(_0859_),
    .X(_0022_));
 sky130_fd_sc_hd__buf_2 _2182_ (.A(_0863_),
    .X(_1322_));
 sky130_fd_sc_hd__nor2_1 _2183_ (.A(_1188_),
    .B(_0886_),
    .Y(_1323_));
 sky130_fd_sc_hd__nor2_4 _2184_ (.A(_0768_),
    .B(_0886_),
    .Y(_1324_));
 sky130_fd_sc_hd__a21oi_4 _2185_ (.A1(_0735_),
    .A2(_0719_),
    .B1(_0737_),
    .Y(_1325_));
 sky130_fd_sc_hd__a21oi_2 _2186_ (.A1(_0854_),
    .A2(_1325_),
    .B1(_0975_),
    .Y(_1326_));
 sky130_fd_sc_hd__or3_1 _2187_ (.A(_1049_),
    .B(_1324_),
    .C(_1326_),
    .X(_1327_));
 sky130_fd_sc_hd__o311a_1 _2188_ (.A1(_1261_),
    .A2(_1202_),
    .A3(_1323_),
    .B1(_1327_),
    .C1(_1178_),
    .X(_1328_));
 sky130_fd_sc_hd__nand2_2 _2189_ (.A(_0918_),
    .B(_0903_),
    .Y(_1329_));
 sky130_fd_sc_hd__nor2_2 _2190_ (.A(_1041_),
    .B(_0976_),
    .Y(_1330_));
 sky130_fd_sc_hd__nor2_1 _2191_ (.A(_1056_),
    .B(_1330_),
    .Y(_1331_));
 sky130_fd_sc_hd__a221o_1 _2192_ (.A1(_0789_),
    .A2(_0876_),
    .B1(_1329_),
    .B2(_1331_),
    .C1(_0915_),
    .X(_1332_));
 sky130_fd_sc_hd__and3b_1 _2193_ (.A_N(_1328_),
    .B(_1164_),
    .C(_1332_),
    .X(_1333_));
 sky130_fd_sc_hd__and3_2 _2194_ (.A(_0763_),
    .B(_0891_),
    .C(_0927_),
    .X(_1334_));
 sky130_fd_sc_hd__clkbuf_4 _2195_ (.A(_1211_),
    .X(_1335_));
 sky130_fd_sc_hd__o21a_1 _2196_ (.A1(_1182_),
    .A2(_1334_),
    .B1(_1335_),
    .X(_1336_));
 sky130_fd_sc_hd__nand2_1 _2197_ (.A(_1291_),
    .B(_0722_),
    .Y(_1337_));
 sky130_fd_sc_hd__o21ai_1 _2198_ (.A1(_1042_),
    .A2(_1337_),
    .B1(_0935_),
    .Y(_1338_));
 sky130_fd_sc_hd__or3_1 _2199_ (.A(_0800_),
    .B(_0890_),
    .C(_1118_),
    .X(_1339_));
 sky130_fd_sc_hd__o32a_2 _2200_ (.A1(_1165_),
    .A2(_0938_),
    .A3(_1141_),
    .B1(_1339_),
    .B2(_1127_),
    .X(_1340_));
 sky130_fd_sc_hd__o221a_1 _2201_ (.A1(_1336_),
    .A2(_1338_),
    .B1(_1340_),
    .B2(_1250_),
    .C1(_0843_),
    .X(_1341_));
 sky130_fd_sc_hd__buf_4 _2202_ (.A(_1115_),
    .X(_1342_));
 sky130_fd_sc_hd__clkbuf_4 _2203_ (.A(_0878_),
    .X(_1343_));
 sky130_fd_sc_hd__nand2_1 _2204_ (.A(_0867_),
    .B(_1030_),
    .Y(_1344_));
 sky130_fd_sc_hd__clkbuf_4 _2205_ (.A(_0936_),
    .X(_1345_));
 sky130_fd_sc_hd__o211a_1 _2206_ (.A1(_1343_),
    .A2(_0868_),
    .B1(_1344_),
    .C1(_1345_),
    .X(_1346_));
 sky130_fd_sc_hd__buf_4 _2207_ (.A(_0786_),
    .X(_1347_));
 sky130_fd_sc_hd__clkbuf_4 _2208_ (.A(_1056_),
    .X(_1348_));
 sky130_fd_sc_hd__o221a_1 _2209_ (.A1(_1088_),
    .A2(_1110_),
    .B1(_1236_),
    .B2(_1347_),
    .C1(_1348_),
    .X(_1349_));
 sky130_fd_sc_hd__nand2_2 _2210_ (.A(_1136_),
    .B(_1173_),
    .Y(_1350_));
 sky130_fd_sc_hd__o2111a_1 _2211_ (.A1(_1199_),
    .A2(_1088_),
    .B1(_0879_),
    .C1(_0882_),
    .D1(_0725_),
    .X(_1351_));
 sky130_fd_sc_hd__a311o_1 _2212_ (.A1(_0734_),
    .A2(_1146_),
    .A3(_1350_),
    .B1(_1351_),
    .C1(_1178_),
    .X(_1352_));
 sky130_fd_sc_hd__o311a_1 _2213_ (.A1(_1342_),
    .A2(_1346_),
    .A3(_1349_),
    .B1(_1352_),
    .C1(_0673_),
    .X(_1353_));
 sky130_fd_sc_hd__and3_4 _2214_ (.A(_0926_),
    .B(_0790_),
    .C(_0947_),
    .X(_1354_));
 sky130_fd_sc_hd__a211o_1 _2215_ (.A1(_0971_),
    .A2(_1079_),
    .B1(_1330_),
    .C1(_0911_),
    .X(_1355_));
 sky130_fd_sc_hd__clkbuf_4 _2216_ (.A(_0782_),
    .X(_1356_));
 sky130_fd_sc_hd__o311ai_1 _2217_ (.A1(_0752_),
    .A2(_1190_),
    .A3(_1354_),
    .B1(_1355_),
    .C1(_1356_),
    .Y(_1357_));
 sky130_fd_sc_hd__a21o_1 _2218_ (.A1(_1123_),
    .A2(_0797_),
    .B1(_0785_),
    .X(_1358_));
 sky130_fd_sc_hd__or3_1 _2219_ (.A(_0737_),
    .B(_1041_),
    .C(_0743_),
    .X(_1359_));
 sky130_fd_sc_hd__nand2_1 _2220_ (.A(_1003_),
    .B(_0770_),
    .Y(_1360_));
 sky130_fd_sc_hd__a21oi_1 _2221_ (.A1(_0919_),
    .A2(_1360_),
    .B1(_1261_),
    .Y(_1361_));
 sky130_fd_sc_hd__a311o_1 _2222_ (.A1(_1274_),
    .A2(_1358_),
    .A3(_1359_),
    .B1(_1361_),
    .C1(_1178_),
    .X(_1362_));
 sky130_fd_sc_hd__a31o_1 _2223_ (.A1(_1273_),
    .A2(_1357_),
    .A3(_1362_),
    .B1(_0645_),
    .X(_1363_));
 sky130_fd_sc_hd__o32a_1 _2224_ (.A1(_0861_),
    .A2(_1333_),
    .A3(_1341_),
    .B1(_1353_),
    .B2(_1363_),
    .X(_1364_));
 sky130_fd_sc_hd__buf_4 _2225_ (.A(_1039_),
    .X(_1365_));
 sky130_fd_sc_hd__nor2_1 _2226_ (.A(_1064_),
    .B(_1275_),
    .Y(_1366_));
 sky130_fd_sc_hd__buf_4 _2227_ (.A(_0975_),
    .X(_1367_));
 sky130_fd_sc_hd__a221o_1 _2228_ (.A1(_1019_),
    .A2(_1072_),
    .B1(_0965_),
    .B2(_1367_),
    .C1(_0751_),
    .X(_1368_));
 sky130_fd_sc_hd__o311a_1 _2229_ (.A1(_1183_),
    .A2(_1299_),
    .A3(_1366_),
    .B1(_1368_),
    .C1(_1308_),
    .X(_1369_));
 sky130_fd_sc_hd__or3_1 _2230_ (.A(_0945_),
    .B(_0733_),
    .C(_1305_),
    .X(_1370_));
 sky130_fd_sc_hd__o311a_1 _2231_ (.A1(_0752_),
    .A2(_1182_),
    .A3(_1277_),
    .B1(_1370_),
    .C1(_1356_),
    .X(_1371_));
 sky130_fd_sc_hd__a211o_1 _2232_ (.A1(_0917_),
    .A2(_1066_),
    .B1(_0940_),
    .C1(_1165_),
    .X(_1372_));
 sky130_fd_sc_hd__or3_1 _2233_ (.A(_1180_),
    .B(_0988_),
    .C(_1200_),
    .X(_1373_));
 sky130_fd_sc_hd__a221o_1 _2234_ (.A1(_1229_),
    .A2(_0965_),
    .B1(_1059_),
    .B2(net56),
    .C1(_1140_),
    .X(_1374_));
 sky130_fd_sc_hd__a221o_1 _2235_ (.A1(_1124_),
    .A2(_1221_),
    .B1(_1097_),
    .B2(_0878_),
    .C1(_0922_),
    .X(_1375_));
 sky130_fd_sc_hd__a31o_1 _2236_ (.A1(_1047_),
    .A2(_1374_),
    .A3(_1375_),
    .B1(_0993_),
    .X(_1376_));
 sky130_fd_sc_hd__a31o_2 _2237_ (.A1(_0783_),
    .A2(_1372_),
    .A3(_1373_),
    .B1(_1376_),
    .X(_1377_));
 sky130_fd_sc_hd__o31a_1 _2238_ (.A1(_1243_),
    .A2(_1369_),
    .A3(_1371_),
    .B1(_1377_),
    .X(_1378_));
 sky130_fd_sc_hd__buf_4 _2239_ (.A(_1077_),
    .X(_1379_));
 sky130_fd_sc_hd__and3_2 _2240_ (.A(_0758_),
    .B(_0831_),
    .C(_0947_),
    .X(_1380_));
 sky130_fd_sc_hd__a211o_1 _2241_ (.A1(_0892_),
    .A2(_1379_),
    .B1(_1380_),
    .C1(_1161_),
    .X(_1381_));
 sky130_fd_sc_hd__o211ai_1 _2242_ (.A1(_1365_),
    .A2(_1378_),
    .B1(_1381_),
    .C1(_1322_),
    .Y(_1382_));
 sky130_fd_sc_hd__o211a_1 _2243_ (.A1(_1322_),
    .A2(_1364_),
    .B1(_1382_),
    .C1(_1242_),
    .X(_0023_));
 sky130_fd_sc_hd__a21o_1 _2244_ (.A1(_0817_),
    .A2(_1379_),
    .B1(_0913_),
    .X(_1383_));
 sky130_fd_sc_hd__or3b_1 _2245_ (.A(_1049_),
    .B(_1050_),
    .C_N(_1350_),
    .X(_1384_));
 sky130_fd_sc_hd__o31a_1 _2246_ (.A1(_0811_),
    .A2(_0966_),
    .A3(_1172_),
    .B1(_1384_),
    .X(_1385_));
 sky130_fd_sc_hd__nor2_1 _2247_ (.A(_1250_),
    .B(_1385_),
    .Y(_1386_));
 sky130_fd_sc_hd__a211o_1 _2248_ (.A1(_1229_),
    .A2(_0965_),
    .B1(_1230_),
    .C1(_0923_),
    .X(_1387_));
 sky130_fd_sc_hd__o311a_1 _2249_ (.A1(_1244_),
    .A2(_1326_),
    .A3(_1323_),
    .B1(_1387_),
    .C1(_1356_),
    .X(_1388_));
 sky130_fd_sc_hd__a21o_1 _2250_ (.A1(_0786_),
    .A2(_1031_),
    .B1(_0875_),
    .X(_1389_));
 sky130_fd_sc_hd__a311o_1 _2251_ (.A1(_0892_),
    .A2(_0973_),
    .A3(_1324_),
    .B1(_1267_),
    .C1(_1040_),
    .X(_1390_));
 sky130_fd_sc_hd__nor2_4 _2252_ (.A(_0729_),
    .B(_0730_),
    .Y(_1391_));
 sky130_fd_sc_hd__or3_4 _2253_ (.A(_0726_),
    .B(_1391_),
    .C(_1031_),
    .X(_1392_));
 sky130_fd_sc_hd__a21o_1 _2254_ (.A1(_1020_),
    .A2(_1392_),
    .B1(_1083_),
    .X(_1393_));
 sky130_fd_sc_hd__o211a_1 _2255_ (.A1(_1175_),
    .A2(_1225_),
    .B1(_1393_),
    .C1(_0963_),
    .X(_1394_));
 sky130_fd_sc_hd__a311o_1 _2256_ (.A1(_1285_),
    .A2(_1389_),
    .A3(_1390_),
    .B1(_1394_),
    .C1(_1318_),
    .X(_1395_));
 sky130_fd_sc_hd__clkbuf_4 _2257_ (.A(_1036_),
    .X(_1396_));
 sky130_fd_sc_hd__o311a_1 _2258_ (.A1(_1298_),
    .A2(_1386_),
    .A3(_1388_),
    .B1(_1395_),
    .C1(_1396_),
    .X(_1397_));
 sky130_fd_sc_hd__a21oi_1 _2259_ (.A1(_1365_),
    .A2(_1383_),
    .B1(_1397_),
    .Y(_1398_));
 sky130_fd_sc_hd__nand2_8 _2260_ (.A(_0741_),
    .B(_0996_),
    .Y(_1399_));
 sky130_fd_sc_hd__nor2_1 _2261_ (.A(_1011_),
    .B(_1399_),
    .Y(_1400_));
 sky130_fd_sc_hd__nand2_1 _2262_ (.A(_0802_),
    .B(_1105_),
    .Y(_1401_));
 sky130_fd_sc_hd__and2b_1 _2263_ (.A_N(_1189_),
    .B(_1401_),
    .X(_1402_));
 sky130_fd_sc_hd__buf_4 _2264_ (.A(_1180_),
    .X(_1403_));
 sky130_fd_sc_hd__o221a_1 _2265_ (.A1(_0889_),
    .A2(_1400_),
    .B1(_1402_),
    .B2(_1403_),
    .C1(_0935_),
    .X(_1404_));
 sky130_fd_sc_hd__a211o_1 _2266_ (.A1(_1232_),
    .A2(_1311_),
    .B1(_0787_),
    .C1(_0801_),
    .X(_1405_));
 sky130_fd_sc_hd__o211a_1 _2267_ (.A1(_1244_),
    .A2(_1181_),
    .B1(_1405_),
    .C1(_1310_),
    .X(_1406_));
 sky130_fd_sc_hd__and3_4 _2268_ (.A(_0718_),
    .B(_0763_),
    .C(_0732_),
    .X(_1407_));
 sky130_fd_sc_hd__a211o_1 _2269_ (.A1(_1367_),
    .A2(_1025_),
    .B1(_1407_),
    .C1(_1040_),
    .X(_1408_));
 sky130_fd_sc_hd__a211o_1 _2270_ (.A1(_1073_),
    .A2(_1379_),
    .B1(_1180_),
    .C1(_1066_),
    .X(_1409_));
 sky130_fd_sc_hd__nor2_4 _2271_ (.A(_1015_),
    .B(_0961_),
    .Y(_1410_));
 sky130_fd_sc_hd__a211o_1 _2272_ (.A1(_1011_),
    .A2(_1097_),
    .B1(_1301_),
    .C1(_0750_),
    .X(_1411_));
 sky130_fd_sc_hd__o311a_1 _2273_ (.A1(_0945_),
    .A2(_1119_),
    .A3(_1410_),
    .B1(_1411_),
    .C1(_0963_),
    .X(_1412_));
 sky130_fd_sc_hd__a311o_1 _2274_ (.A1(_0779_),
    .A2(_1408_),
    .A3(_1409_),
    .B1(_1412_),
    .C1(_0667_),
    .X(_1413_));
 sky130_fd_sc_hd__o311a_1 _2275_ (.A1(_1298_),
    .A2(_1404_),
    .A3(_1406_),
    .B1(_1413_),
    .C1(_1396_),
    .X(_1414_));
 sky130_fd_sc_hd__a211o_1 _2276_ (.A1(_0917_),
    .A2(_0816_),
    .B1(_1042_),
    .C1(_1264_),
    .X(_1415_));
 sky130_fd_sc_hd__o311a_1 _2277_ (.A1(_1348_),
    .A2(_0925_),
    .A3(_1380_),
    .B1(_1415_),
    .C1(_1310_),
    .X(_1416_));
 sky130_fd_sc_hd__and3_1 _2278_ (.A(_1367_),
    .B(_0803_),
    .C(_0819_),
    .X(_1417_));
 sky130_fd_sc_hd__and3_1 _2279_ (.A(_0881_),
    .B(_0918_),
    .C(_0797_),
    .X(_1418_));
 sky130_fd_sc_hd__a211o_1 _2280_ (.A1(_1078_),
    .A2(_1229_),
    .B1(_1418_),
    .C1(_0801_),
    .X(_1419_));
 sky130_fd_sc_hd__o311a_1 _2281_ (.A1(_1281_),
    .A2(_1247_),
    .A3(_1417_),
    .B1(_1419_),
    .C1(_1356_),
    .X(_1420_));
 sky130_fd_sc_hd__a221o_1 _2282_ (.A1(_0739_),
    .A2(_0744_),
    .B1(_0816_),
    .B2(_1078_),
    .C1(_0923_),
    .X(_1421_));
 sky130_fd_sc_hd__nor3_4 _2283_ (.A(_0728_),
    .B(_0720_),
    .C(_1007_),
    .Y(_1422_));
 sky130_fd_sc_hd__a221o_1 _2284_ (.A1(_0452_),
    .A2(_0813_),
    .B1(net51),
    .B2(_1232_),
    .C1(_1165_),
    .X(_1423_));
 sky130_fd_sc_hd__a211o_1 _2285_ (.A1(_1000_),
    .A2(_1229_),
    .B1(_1176_),
    .C1(_1140_),
    .X(_1424_));
 sky130_fd_sc_hd__a211o_1 _2286_ (.A1(_0947_),
    .A2(_0948_),
    .B1(_1314_),
    .C1(_1083_),
    .X(_1425_));
 sky130_fd_sc_hd__a31o_1 _2287_ (.A1(_1047_),
    .A2(_1424_),
    .A3(_1425_),
    .B1(_0842_),
    .X(_1426_));
 sky130_fd_sc_hd__a31o_1 _2288_ (.A1(_0783_),
    .A2(_1421_),
    .A3(_1423_),
    .B1(_1426_),
    .X(_1427_));
 sky130_fd_sc_hd__o311a_1 _2289_ (.A1(_0673_),
    .A2(_1416_),
    .A3(_1420_),
    .B1(_1427_),
    .C1(_0861_),
    .X(_1428_));
 sky130_fd_sc_hd__o21ai_1 _2290_ (.A1(_1414_),
    .A2(_1428_),
    .B1(_1197_),
    .Y(_1429_));
 sky130_fd_sc_hd__o211a_1 _2291_ (.A1(_1158_),
    .A2(_1398_),
    .B1(_1429_),
    .C1(_1242_),
    .X(_0024_));
 sky130_fd_sc_hd__a21o_1 _2292_ (.A1(_1067_),
    .A2(_1401_),
    .B1(_0754_),
    .X(_1430_));
 sky130_fd_sc_hd__o311a_1 _2293_ (.A1(_0985_),
    .A2(_1200_),
    .A3(_1302_),
    .B1(_1430_),
    .C1(_0777_),
    .X(_1431_));
 sky130_fd_sc_hd__and3_4 _2294_ (.A(_0728_),
    .B(_1078_),
    .C(_0996_),
    .X(_1432_));
 sky130_fd_sc_hd__and3_1 _2295_ (.A(_0772_),
    .B(_0926_),
    .C(_1391_),
    .X(_1433_));
 sky130_fd_sc_hd__or3b_1 _2296_ (.A(_1305_),
    .B(_0749_),
    .C_N(_0961_),
    .X(_1434_));
 sky130_fd_sc_hd__o311a_1 _2297_ (.A1(_1140_),
    .A2(_1432_),
    .A3(_1433_),
    .B1(_1434_),
    .C1(_0694_),
    .X(_1435_));
 sky130_fd_sc_hd__a221o_1 _2298_ (.A1(_0806_),
    .A2(_1020_),
    .B1(_1097_),
    .B2(_1117_),
    .C1(_0835_),
    .X(_1436_));
 sky130_fd_sc_hd__o311a_1 _2299_ (.A1(_0810_),
    .A2(_1103_),
    .A3(_1302_),
    .B1(_1436_),
    .C1(_0694_),
    .X(_1437_));
 sky130_fd_sc_hd__nor2_1 _2300_ (.A(_0877_),
    .B(_0903_),
    .Y(_1438_));
 sky130_fd_sc_hd__and3_1 _2301_ (.A(_0716_),
    .B(_0829_),
    .C(net56),
    .X(_1439_));
 sky130_fd_sc_hd__o32a_1 _2302_ (.A1(_0964_),
    .A2(_1438_),
    .A3(_1439_),
    .B1(_1292_),
    .B2(_0900_),
    .X(_1440_));
 sky130_fd_sc_hd__o21ai_1 _2303_ (.A1(_0963_),
    .A2(_1440_),
    .B1(_0993_),
    .Y(_1441_));
 sky130_fd_sc_hd__o32a_1 _2304_ (.A1(_0993_),
    .A2(_1431_),
    .A3(_1435_),
    .B1(_1437_),
    .B2(_1441_),
    .X(_1442_));
 sky130_fd_sc_hd__and3_2 _2305_ (.A(_1003_),
    .B(_0939_),
    .C(_0790_),
    .X(_1443_));
 sky130_fd_sc_hd__a31o_1 _2306_ (.A1(_1089_),
    .A2(_1343_),
    .A3(_0929_),
    .B1(_1443_),
    .X(_1444_));
 sky130_fd_sc_hd__or4_1 _2307_ (.A(_0835_),
    .B(_1249_),
    .C(_1050_),
    .D(_1410_),
    .X(_1445_));
 sky130_fd_sc_hd__a311o_1 _2308_ (.A1(_1003_),
    .A2(_0878_),
    .A3(_1013_),
    .B1(_1294_),
    .C1(_0922_),
    .X(_1446_));
 sky130_fd_sc_hd__a21oi_1 _2309_ (.A1(_1445_),
    .A2(_1446_),
    .B1(_0915_),
    .Y(_1447_));
 sky130_fd_sc_hd__nor2_2 _2310_ (.A(_1117_),
    .B(_1097_),
    .Y(_1448_));
 sky130_fd_sc_hd__nor2_2 _2311_ (.A(_1052_),
    .B(_1167_),
    .Y(_1449_));
 sky130_fd_sc_hd__o21ai_1 _2312_ (.A1(_1448_),
    .A2(_1449_),
    .B1(_1235_),
    .Y(_1450_));
 sky130_fd_sc_hd__or3b_1 _2313_ (.A(_0835_),
    .B(_1249_),
    .C_N(_1085_),
    .X(_1451_));
 sky130_fd_sc_hd__a31o_1 _2314_ (.A1(_0934_),
    .A2(_1450_),
    .A3(_1451_),
    .B1(_0841_),
    .X(_1452_));
 sky130_fd_sc_hd__nand2_1 _2315_ (.A(_0721_),
    .B(_0829_),
    .Y(_1453_));
 sky130_fd_sc_hd__o221a_1 _2316_ (.A1(_0787_),
    .A2(_1188_),
    .B1(_0869_),
    .B2(_1236_),
    .C1(_0984_),
    .X(_1454_));
 sky130_fd_sc_hd__a31o_1 _2317_ (.A1(_0800_),
    .A2(_1001_),
    .A3(_1453_),
    .B1(_1454_),
    .X(_1455_));
 sky130_fd_sc_hd__nor2_1 _2318_ (.A(_0743_),
    .B(_1001_),
    .Y(_1456_));
 sky130_fd_sc_hd__and3_2 _2319_ (.A(_0852_),
    .B(_0727_),
    .C(_0996_),
    .X(_1457_));
 sky130_fd_sc_hd__or3_1 _2320_ (.A(_0723_),
    .B(_1066_),
    .C(_1457_),
    .X(_1458_));
 sky130_fd_sc_hd__o311a_1 _2321_ (.A1(_0910_),
    .A2(_1175_),
    .A3(_1456_),
    .B1(_1458_),
    .C1(_0685_),
    .X(_1459_));
 sky130_fd_sc_hd__a211o_1 _2322_ (.A1(_0934_),
    .A2(_1455_),
    .B1(_1459_),
    .C1(_0661_),
    .X(_1460_));
 sky130_fd_sc_hd__o21ai_1 _2323_ (.A1(_1447_),
    .A2(_1452_),
    .B1(_1460_),
    .Y(_1461_));
 sky130_fd_sc_hd__a21oi_2 _2324_ (.A1(_0854_),
    .A2(_1325_),
    .B1(_1041_),
    .Y(_1462_));
 sky130_fd_sc_hd__nor2_1 _2325_ (.A(_0791_),
    .B(_0805_),
    .Y(_1463_));
 sky130_fd_sc_hd__a211o_1 _2326_ (.A1(_1123_),
    .A2(_1106_),
    .B1(_1463_),
    .C1(_0799_),
    .X(_1464_));
 sky130_fd_sc_hd__o311a_1 _2327_ (.A1(_0985_),
    .A2(_1407_),
    .A3(_1462_),
    .B1(_1464_),
    .C1(_0838_),
    .X(_1465_));
 sky130_fd_sc_hd__and2b_4 _2328_ (.A_N(_1159_),
    .B(_1032_),
    .X(_1466_));
 sky130_fd_sc_hd__and3_2 _2329_ (.A(_0772_),
    .B(_0758_),
    .C(_0790_),
    .X(_1467_));
 sky130_fd_sc_hd__or3_1 _2330_ (.A(_0834_),
    .B(_0888_),
    .C(_1301_),
    .X(_1468_));
 sky130_fd_sc_hd__o311a_1 _2331_ (.A1(_0922_),
    .A2(_1466_),
    .A3(_1467_),
    .B1(_1468_),
    .C1(_0914_),
    .X(_1469_));
 sky130_fd_sc_hd__and3_2 _2332_ (.A(_0740_),
    .B(_0854_),
    .C(_0897_),
    .X(_1470_));
 sky130_fd_sc_hd__a211o_1 _2333_ (.A1(_1013_),
    .A2(_1205_),
    .B1(_1470_),
    .C1(_0754_),
    .X(_1471_));
 sky130_fd_sc_hd__a221o_1 _2334_ (.A1(_0828_),
    .A2(_1084_),
    .B1(_1127_),
    .B2(_0823_),
    .C1(_0864_),
    .X(_1472_));
 sky130_fd_sc_hd__and3_1 _2335_ (.A(_0694_),
    .B(_1471_),
    .C(_1472_),
    .X(_1473_));
 sky130_fd_sc_hd__a211o_1 _2336_ (.A1(_0797_),
    .A2(_1084_),
    .B1(_1150_),
    .C1(_0835_),
    .X(_1474_));
 sky130_fd_sc_hd__nor2_4 _2337_ (.A(_0728_),
    .B(_1391_),
    .Y(_1475_));
 sky130_fd_sc_hd__or3b_1 _2338_ (.A(_0799_),
    .B(_1475_),
    .C_N(_1054_),
    .X(_1476_));
 sky130_fd_sc_hd__a31o_1 _2339_ (.A1(_0914_),
    .A2(_1474_),
    .A3(_1476_),
    .B1(_0661_),
    .X(_1477_));
 sky130_fd_sc_hd__o32a_1 _2340_ (.A1(_0842_),
    .A2(_1465_),
    .A3(_1469_),
    .B1(_1473_),
    .B2(_1477_),
    .X(_1478_));
 sky130_fd_sc_hd__mux4_1 _2341_ (.A0(_1442_),
    .A1(_1444_),
    .A2(_1461_),
    .A3(_1478_),
    .S0(_0863_),
    .S1(_0645_),
    .X(_1479_));
 sky130_fd_sc_hd__and2b_1 _2342_ (.A_N(_1479_),
    .B(_0859_),
    .X(_1480_));
 sky130_fd_sc_hd__clkbuf_1 _2343_ (.A(_1480_),
    .X(_0025_));
 sky130_fd_sc_hd__o21ai_1 _2344_ (.A1(_1347_),
    .A2(_1088_),
    .B1(_1054_),
    .Y(_1481_));
 sky130_fd_sc_hd__or3_2 _2345_ (.A(_0911_),
    .B(_0774_),
    .C(_1467_),
    .X(_1482_));
 sky130_fd_sc_hd__a21o_1 _2346_ (.A1(_1160_),
    .A2(_1344_),
    .B1(_1291_),
    .X(_1483_));
 sky130_fd_sc_hd__a21oi_1 _2347_ (.A1(_1482_),
    .A2(_1483_),
    .B1(_1342_),
    .Y(_1484_));
 sky130_fd_sc_hd__a211o_1 _2348_ (.A1(_1073_),
    .A2(_1379_),
    .B1(_1439_),
    .C1(_0923_),
    .X(_1485_));
 sky130_fd_sc_hd__o311a_1 _2349_ (.A1(_1244_),
    .A2(_0733_),
    .A3(_0813_),
    .B1(_1485_),
    .C1(_1342_),
    .X(_1486_));
 sky130_fd_sc_hd__and3_1 _2350_ (.A(_0825_),
    .B(_0820_),
    .C(_1025_),
    .X(_1487_));
 sky130_fd_sc_hd__or4_1 _2351_ (.A(_0810_),
    .B(_1050_),
    .C(_1410_),
    .D(_1487_),
    .X(_1488_));
 sky130_fd_sc_hd__a211o_1 _2352_ (.A1(_0816_),
    .A2(_0817_),
    .B1(_1448_),
    .C1(_1264_),
    .X(_1489_));
 sky130_fd_sc_hd__nor2_1 _2353_ (.A(_1078_),
    .B(_1059_),
    .Y(_1490_));
 sky130_fd_sc_hd__nor2_4 _2354_ (.A(_0728_),
    .B(_0829_),
    .Y(_1491_));
 sky130_fd_sc_hd__a211o_1 _2355_ (.A1(_1000_),
    .A2(_1043_),
    .B1(_1491_),
    .C1(_0800_),
    .X(_1492_));
 sky130_fd_sc_hd__o311a_1 _2356_ (.A1(_0945_),
    .A2(_1002_),
    .A3(_1490_),
    .B1(_1492_),
    .C1(_0978_),
    .X(_1493_));
 sky130_fd_sc_hd__a311o_4 _2357_ (.A1(_1308_),
    .A2(_1488_),
    .A3(_1489_),
    .B1(_1493_),
    .C1(_1318_),
    .X(_1494_));
 sky130_fd_sc_hd__o311a_1 _2358_ (.A1(_1298_),
    .A2(_1484_),
    .A3(_1486_),
    .B1(_1494_),
    .C1(_1396_),
    .X(_1495_));
 sky130_fd_sc_hd__a21oi_1 _2359_ (.A1(_1365_),
    .A2(_1481_),
    .B1(_1495_),
    .Y(_1496_));
 sky130_fd_sc_hd__or2_2 _2360_ (.A(_0769_),
    .B(_1073_),
    .X(_1497_));
 sky130_fd_sc_hd__nand3_1 _2361_ (.A(_1335_),
    .B(_1107_),
    .C(_1497_),
    .Y(_1498_));
 sky130_fd_sc_hd__o311a_1 _2362_ (.A1(_1345_),
    .A2(_0898_),
    .A3(_0948_),
    .B1(_1498_),
    .C1(_1287_),
    .X(_1499_));
 sky130_fd_sc_hd__and3_2 _2363_ (.A(_1089_),
    .B(_0713_),
    .C(_0744_),
    .X(_1500_));
 sky130_fd_sc_hd__nor2_1 _2364_ (.A(_0770_),
    .B(_0788_),
    .Y(_1501_));
 sky130_fd_sc_hd__or3_1 _2365_ (.A(_0936_),
    .B(_0988_),
    .C(_1200_),
    .X(_1502_));
 sky130_fd_sc_hd__o311a_1 _2366_ (.A1(_1403_),
    .A2(_1500_),
    .A3(_1501_),
    .B1(_0935_),
    .C1(_1502_),
    .X(_1503_));
 sky130_fd_sc_hd__a221o_1 _2367_ (.A1(_1311_),
    .A2(_0867_),
    .B1(_0892_),
    .B2(_1379_),
    .C1(_1180_),
    .X(_1504_));
 sky130_fd_sc_hd__a211o_1 _2368_ (.A1(_1311_),
    .A2(net52),
    .B1(_1026_),
    .C1(_1040_),
    .X(_1505_));
 sky130_fd_sc_hd__nand2_1 _2369_ (.A(_0892_),
    .B(_0973_),
    .Y(_1506_));
 sky130_fd_sc_hd__a221o_1 _2370_ (.A1(_0916_),
    .A2(_0815_),
    .B1(_1506_),
    .B2(_0970_),
    .C1(_1028_),
    .X(_1507_));
 sky130_fd_sc_hd__o311a_1 _2371_ (.A1(_0957_),
    .A2(_1283_),
    .A3(_1448_),
    .B1(_1507_),
    .C1(_0963_),
    .X(_1508_));
 sky130_fd_sc_hd__a311o_1 _2372_ (.A1(_0779_),
    .A2(_1504_),
    .A3(_1505_),
    .B1(_1508_),
    .C1(_0667_),
    .X(_1509_));
 sky130_fd_sc_hd__o311a_1 _2373_ (.A1(_1273_),
    .A2(_1499_),
    .A3(_1503_),
    .B1(_1509_),
    .C1(_1396_),
    .X(_1510_));
 sky130_fd_sc_hd__and2_1 _2374_ (.A(_1117_),
    .B(net52),
    .X(_1511_));
 sky130_fd_sc_hd__nor2_1 _2375_ (.A(_1078_),
    .B(_1392_),
    .Y(_1512_));
 sky130_fd_sc_hd__or3b_1 _2376_ (.A(_1512_),
    .B(_0725_),
    .C_N(_0761_),
    .X(_1513_));
 sky130_fd_sc_hd__o311a_1 _2377_ (.A1(_1281_),
    .A2(_1491_),
    .A3(_1511_),
    .B1(_1513_),
    .C1(_1310_),
    .X(_1514_));
 sky130_fd_sc_hd__a211o_1 _2378_ (.A1(_1012_),
    .A2(_1347_),
    .B1(_1202_),
    .C1(_1291_),
    .X(_1515_));
 sky130_fd_sc_hd__and3_1 _2379_ (.A(_0975_),
    .B(_0924_),
    .C(_0851_),
    .X(_1516_));
 sky130_fd_sc_hd__or3_1 _2380_ (.A(_0911_),
    .B(_0990_),
    .C(_1516_),
    .X(_1517_));
 sky130_fd_sc_hd__a21oi_1 _2381_ (.A1(_1515_),
    .A2(_1517_),
    .B1(_0706_),
    .Y(_1518_));
 sky130_fd_sc_hd__nand2_1 _2382_ (.A(_0807_),
    .B(_0976_),
    .Y(_1519_));
 sky130_fd_sc_hd__nand2_1 _2383_ (.A(_1043_),
    .B(_0916_),
    .Y(_1520_));
 sky130_fd_sc_hd__nand3_1 _2384_ (.A(_1335_),
    .B(_1519_),
    .C(_1520_),
    .Y(_1521_));
 sky130_fd_sc_hd__a221o_1 _2385_ (.A1(_0803_),
    .A2(_0816_),
    .B1(_1030_),
    .B2(_0735_),
    .C1(_1040_),
    .X(_1522_));
 sky130_fd_sc_hd__and3_1 _2386_ (.A(_0852_),
    .B(_0970_),
    .C(_1025_),
    .X(_1523_));
 sky130_fd_sc_hd__and3_2 _2387_ (.A(_1015_),
    .B(_0823_),
    .C(_0738_),
    .X(_1524_));
 sky130_fd_sc_hd__a211o_1 _2388_ (.A1(_0806_),
    .A2(_1020_),
    .B1(_1524_),
    .C1(_1060_),
    .X(_1525_));
 sky130_fd_sc_hd__o311a_1 _2389_ (.A1(_0957_),
    .A2(_1043_),
    .A3(_1523_),
    .B1(_1525_),
    .C1(_0978_),
    .X(_1526_));
 sky130_fd_sc_hd__a311o_1 _2390_ (.A1(_1310_),
    .A2(_1521_),
    .A3(_1522_),
    .B1(_1526_),
    .C1(_1318_),
    .X(_1527_));
 sky130_fd_sc_hd__o311a_1 _2391_ (.A1(_1298_),
    .A2(_1514_),
    .A3(_1518_),
    .B1(_1527_),
    .C1(_0861_),
    .X(_1528_));
 sky130_fd_sc_hd__o21ai_1 _2392_ (.A1(_1510_),
    .A2(_1528_),
    .B1(_1197_),
    .Y(_1529_));
 sky130_fd_sc_hd__o211a_1 _2393_ (.A1(_1158_),
    .A2(_1496_),
    .B1(_1529_),
    .C1(_1242_),
    .X(_0026_));
 sky130_fd_sc_hd__and3_1 _2394_ (.A(_0785_),
    .B(_0713_),
    .C(_0959_),
    .X(_1530_));
 sky130_fd_sc_hd__or3_1 _2395_ (.A(_1256_),
    .B(_1233_),
    .C(_1530_),
    .X(_1531_));
 sky130_fd_sc_hd__nand2_1 _2396_ (.A(_0947_),
    .B(_0931_),
    .Y(_1532_));
 sky130_fd_sc_hd__a21o_1 _2397_ (.A1(_1532_),
    .A2(_1350_),
    .B1(_0752_),
    .X(_0059_));
 sky130_fd_sc_hd__a211o_1 _2398_ (.A1(_1003_),
    .A2(_1311_),
    .B1(_1516_),
    .C1(_1109_),
    .X(_0060_));
 sky130_fd_sc_hd__o311a_1 _2399_ (.A1(_1274_),
    .A2(_1042_),
    .A3(_1129_),
    .B1(_0060_),
    .C1(_1278_),
    .X(_0061_));
 sky130_fd_sc_hd__a311o_1 _2400_ (.A1(_1250_),
    .A2(_1531_),
    .A3(_0059_),
    .B1(_0061_),
    .C1(_1273_),
    .X(_0062_));
 sky130_fd_sc_hd__or3b_2 _2401_ (.A(_1276_),
    .B(_0811_),
    .C_N(_1085_),
    .X(_0063_));
 sky130_fd_sc_hd__or3_1 _2402_ (.A(_1256_),
    .B(_0980_),
    .C(_1283_),
    .X(_0064_));
 sky130_fd_sc_hd__o221a_1 _2403_ (.A1(_1225_),
    .A2(_1294_),
    .B1(_1253_),
    .B2(_1400_),
    .C1(_1178_),
    .X(_0065_));
 sky130_fd_sc_hd__a311o_1 _2404_ (.A1(_0706_),
    .A2(_0063_),
    .A3(_0064_),
    .B1(_0065_),
    .C1(_1164_),
    .X(_0066_));
 sky130_fd_sc_hd__a21oi_2 _2405_ (.A1(_0062_),
    .A2(_0066_),
    .B1(_1365_),
    .Y(_0067_));
 sky130_fd_sc_hd__o211a_1 _2406_ (.A1(_1110_),
    .A2(_0886_),
    .B1(_0879_),
    .C1(_1365_),
    .X(_0068_));
 sky130_fd_sc_hd__or3_1 _2407_ (.A(_1391_),
    .B(_0880_),
    .C(_0900_),
    .X(_0069_));
 sky130_fd_sc_hd__a21o_1 _2408_ (.A1(_1110_),
    .A2(_1020_),
    .B1(_0911_),
    .X(_0070_));
 sky130_fd_sc_hd__a211o_1 _2409_ (.A1(_1113_),
    .A2(_1072_),
    .B1(_1150_),
    .C1(_1028_),
    .X(_0071_));
 sky130_fd_sc_hd__a211o_1 _2410_ (.A1(_1089_),
    .A2(_0970_),
    .B1(_0893_),
    .C1(_0750_),
    .X(_0072_));
 sky130_fd_sc_hd__a31o_1 _2411_ (.A1(_0934_),
    .A2(_0071_),
    .A3(_0072_),
    .B1(_0661_),
    .X(_0073_));
 sky130_fd_sc_hd__a31o_1 _2412_ (.A1(_1287_),
    .A2(_0069_),
    .A3(_0070_),
    .B1(_0073_),
    .X(_0074_));
 sky130_fd_sc_hd__nor2_4 _2413_ (.A(_0728_),
    .B(_1181_),
    .Y(_0075_));
 sky130_fd_sc_hd__and3_2 _2414_ (.A(_0765_),
    .B(_0784_),
    .C(_0719_),
    .X(_0076_));
 sky130_fd_sc_hd__or3_1 _2415_ (.A(_0984_),
    .B(_1202_),
    .C(_0076_),
    .X(_0077_));
 sky130_fd_sc_hd__o311a_1 _2416_ (.A1(_0755_),
    .A2(_0832_),
    .A3(_0075_),
    .B1(_0077_),
    .C1(_0694_),
    .X(_0078_));
 sky130_fd_sc_hd__a31o_1 _2417_ (.A1(_0820_),
    .A2(_0738_),
    .A3(_0937_),
    .B1(_1325_),
    .X(_0079_));
 sky130_fd_sc_hd__a31o_2 _2418_ (.A1(_0831_),
    .A2(_0892_),
    .A3(_0973_),
    .B1(_0740_),
    .X(_0080_));
 sky130_fd_sc_hd__and3b_1 _2419_ (.A_N(_1090_),
    .B(_0080_),
    .C(_0984_),
    .X(_0081_));
 sky130_fd_sc_hd__a311o_1 _2420_ (.A1(_0810_),
    .A2(_1160_),
    .A3(_0079_),
    .B1(_0081_),
    .C1(_0838_),
    .X(_0082_));
 sky130_fd_sc_hd__or3b_2 _2421_ (.A(_0842_),
    .B(_0078_),
    .C_N(_0082_),
    .X(_0083_));
 sky130_fd_sc_hd__a21oi_1 _2422_ (.A1(_0074_),
    .A2(_0083_),
    .B1(_1161_),
    .Y(_0084_));
 sky130_fd_sc_hd__and2b_1 _2423_ (.A_N(_1443_),
    .B(_0080_),
    .X(_0085_));
 sky130_fd_sc_hd__a31o_1 _2424_ (.A1(_1011_),
    .A2(_0971_),
    .A3(_0973_),
    .B1(_0750_),
    .X(_0086_));
 sky130_fd_sc_hd__o221a_1 _2425_ (.A1(_1165_),
    .A2(_0085_),
    .B1(_0086_),
    .B2(_0744_),
    .C1(_0839_),
    .X(_0087_));
 sky130_fd_sc_hd__or3b_1 _2426_ (.A(_1235_),
    .B(_0962_),
    .C_N(_1097_),
    .X(_0088_));
 sky130_fd_sc_hd__or3_1 _2427_ (.A(_0810_),
    .B(_1439_),
    .C(_1443_),
    .X(_0089_));
 sky130_fd_sc_hd__a21oi_1 _2428_ (.A1(_0088_),
    .A2(_0089_),
    .B1(_1278_),
    .Y(_0090_));
 sky130_fd_sc_hd__a221o_1 _2429_ (.A1(_0999_),
    .A2(_1221_),
    .B1(_1112_),
    .B2(_1219_),
    .C1(_0910_),
    .X(_0091_));
 sky130_fd_sc_hd__o31ai_1 _2430_ (.A1(_0875_),
    .A2(_1189_),
    .A3(_1380_),
    .B1(_0091_),
    .Y(_0092_));
 sky130_fd_sc_hd__or3_2 _2431_ (.A(_0716_),
    .B(_0896_),
    .C(_1052_),
    .X(_0093_));
 sky130_fd_sc_hd__o221a_1 _2432_ (.A1(_0965_),
    .A2(_1275_),
    .B1(_0093_),
    .B2(_1083_),
    .C1(_0914_),
    .X(_0094_));
 sky130_fd_sc_hd__a221o_1 _2433_ (.A1(_0839_),
    .A2(_0092_),
    .B1(_0094_),
    .B2(_1098_),
    .C1(_0907_),
    .X(_0095_));
 sky130_fd_sc_hd__o311a_1 _2434_ (.A1(_0843_),
    .A2(_0087_),
    .A3(_0090_),
    .B1(_0095_),
    .C1(_0645_),
    .X(_0096_));
 sky130_fd_sc_hd__or3_1 _2435_ (.A(_0863_),
    .B(_0084_),
    .C(_0096_),
    .X(_0097_));
 sky130_fd_sc_hd__o311a_1 _2436_ (.A1(_1158_),
    .A2(_0067_),
    .A3(_0068_),
    .B1(_0859_),
    .C1(_0097_),
    .X(_0027_));
 sky130_fd_sc_hd__nand2_1 _2437_ (.A(_0871_),
    .B(_1360_),
    .Y(_0098_));
 sky130_fd_sc_hd__mux2_1 _2438_ (.A0(_1335_),
    .A1(_1248_),
    .S(_0098_),
    .X(_0099_));
 sky130_fd_sc_hd__or3b_1 _2439_ (.A(_0836_),
    .B(_1045_),
    .C_N(_1497_),
    .X(_0100_));
 sky130_fd_sc_hd__o311a_1 _2440_ (.A1(_1274_),
    .A2(_0733_),
    .A3(_1130_),
    .B1(_0100_),
    .C1(_1198_),
    .X(_0101_));
 sky130_fd_sc_hd__a211o_1 _2441_ (.A1(_0706_),
    .A2(_0099_),
    .B1(_0101_),
    .C1(_1164_),
    .X(_0102_));
 sky130_fd_sc_hd__a31o_1 _2442_ (.A1(_1089_),
    .A2(_1343_),
    .A3(_0929_),
    .B1(_0942_),
    .X(_0103_));
 sky130_fd_sc_hd__a211o_1 _2443_ (.A1(_1343_),
    .A2(_0973_),
    .B1(_0912_),
    .C1(_1335_),
    .X(_0104_));
 sky130_fd_sc_hd__and3_1 _2444_ (.A(_0820_),
    .B(_0829_),
    .C(_1173_),
    .X(_0105_));
 sky130_fd_sc_hd__or3_1 _2445_ (.A(_1049_),
    .B(_1079_),
    .C(_0105_),
    .X(_0106_));
 sky130_fd_sc_hd__o311a_1 _2446_ (.A1(_1291_),
    .A2(net51),
    .A3(_1443_),
    .B1(_0106_),
    .C1(_0703_),
    .X(_0107_));
 sky130_fd_sc_hd__a311o_1 _2447_ (.A1(_1250_),
    .A2(_0103_),
    .A3(_0104_),
    .B1(_0107_),
    .C1(_1273_),
    .X(_0108_));
 sky130_fd_sc_hd__nor2_1 _2448_ (.A(_1120_),
    .B(net56),
    .Y(_0109_));
 sky130_fd_sc_hd__or3_1 _2449_ (.A(_1117_),
    .B(_0813_),
    .C(_0867_),
    .X(_0110_));
 sky130_fd_sc_hd__a21o_1 _2450_ (.A1(_1275_),
    .A2(_0110_),
    .B1(_0751_),
    .X(_0111_));
 sky130_fd_sc_hd__o311a_1 _2451_ (.A1(_1256_),
    .A2(_1282_),
    .A3(_0109_),
    .B1(_0111_),
    .C1(_1278_),
    .X(_0112_));
 sky130_fd_sc_hd__or2_1 _2452_ (.A(_1235_),
    .B(_1294_),
    .X(_0113_));
 sky130_fd_sc_hd__o221a_1 _2453_ (.A1(_1023_),
    .A2(_1253_),
    .B1(_0113_),
    .B2(_1135_),
    .C1(_1198_),
    .X(_0114_));
 sky130_fd_sc_hd__a21o_1 _2454_ (.A1(_1019_),
    .A2(_0855_),
    .B1(_1060_),
    .X(_0115_));
 sky130_fd_sc_hd__a21o_1 _2455_ (.A1(_0086_),
    .A2(_0115_),
    .B1(_0764_),
    .X(_0116_));
 sky130_fd_sc_hd__a221o_1 _2456_ (.A1(_1136_),
    .A2(_0738_),
    .B1(_0929_),
    .B2(_1206_),
    .C1(_0956_),
    .X(_0117_));
 sky130_fd_sc_hd__o311a_1 _2457_ (.A1(_0936_),
    .A2(_0798_),
    .A3(_1112_),
    .B1(_0117_),
    .C1(_0934_),
    .X(_0118_));
 sky130_fd_sc_hd__a211o_1 _2458_ (.A1(_1278_),
    .A2(_0116_),
    .B1(_0118_),
    .C1(_0907_),
    .X(_0119_));
 sky130_fd_sc_hd__o311a_1 _2459_ (.A1(_1273_),
    .A2(_0112_),
    .A3(_0114_),
    .B1(_0119_),
    .C1(_1161_),
    .X(_0120_));
 sky130_fd_sc_hd__a31oi_2 _2460_ (.A1(_1365_),
    .A2(_0102_),
    .A3(_0108_),
    .B1(_0120_),
    .Y(_0121_));
 sky130_fd_sc_hd__or3_1 _2461_ (.A(_0836_),
    .B(_1289_),
    .C(_1462_),
    .X(_0122_));
 sky130_fd_sc_hd__o311a_1 _2462_ (.A1(_1291_),
    .A2(_1448_),
    .A3(_1511_),
    .B1(_0122_),
    .C1(_1198_),
    .X(_0123_));
 sky130_fd_sc_hd__nor2_4 _2463_ (.A(_1011_),
    .B(_0903_),
    .Y(_0124_));
 sky130_fd_sc_hd__or3_1 _2464_ (.A(_1063_),
    .B(_1053_),
    .C(_1277_),
    .X(_0125_));
 sky130_fd_sc_hd__o311a_1 _2465_ (.A1(_1335_),
    .A2(_0124_),
    .A3(_1457_),
    .B1(_0125_),
    .C1(_1278_),
    .X(_0126_));
 sky130_fd_sc_hd__or3_1 _2466_ (.A(_1273_),
    .B(_0123_),
    .C(_0126_),
    .X(_0127_));
 sky130_fd_sc_hd__o21a_1 _2467_ (.A1(_1168_),
    .A2(_0076_),
    .B1(_0911_),
    .X(_0128_));
 sky130_fd_sc_hd__a31o_1 _2468_ (.A1(_0739_),
    .A2(_0817_),
    .A3(_1220_),
    .B1(_0128_),
    .X(_0129_));
 sky130_fd_sc_hd__nor2_1 _2469_ (.A(_0918_),
    .B(_0896_),
    .Y(_0130_));
 sky130_fd_sc_hd__or3_1 _2470_ (.A(_1211_),
    .B(_1418_),
    .C(_0130_),
    .X(_0131_));
 sky130_fd_sc_hd__o311a_1 _2471_ (.A1(_1348_),
    .A2(_0774_),
    .A3(_1059_),
    .B1(_0131_),
    .C1(_0779_),
    .X(_0132_));
 sky130_fd_sc_hd__a211o_1 _2472_ (.A1(_0706_),
    .A2(_0129_),
    .B1(_0132_),
    .C1(_0673_),
    .X(_0133_));
 sky130_fd_sc_hd__a21oi_1 _2473_ (.A1(_0127_),
    .A2(_0133_),
    .B1(_1365_),
    .Y(_0134_));
 sky130_fd_sc_hd__a31o_1 _2474_ (.A1(_0861_),
    .A2(_1065_),
    .A3(_0093_),
    .B1(_0849_),
    .X(_0135_));
 sky130_fd_sc_hd__o221a_1 _2475_ (.A1(_1322_),
    .A2(_0121_),
    .B1(_0134_),
    .B2(_0135_),
    .C1(_0859_),
    .X(_0005_));
 sky130_fd_sc_hd__or3_1 _2476_ (.A(_1036_),
    .B(_0737_),
    .C(_1343_),
    .X(_0136_));
 sky130_fd_sc_hd__and3_4 _2477_ (.A(_0757_),
    .B(_0712_),
    .C(_0965_),
    .X(_0137_));
 sky130_fd_sc_hd__or3_1 _2478_ (.A(_0956_),
    .B(_1094_),
    .C(_0137_),
    .X(_0138_));
 sky130_fd_sc_hd__o31a_1 _2479_ (.A1(_1264_),
    .A2(_1111_),
    .A3(_1500_),
    .B1(_0138_),
    .X(_0139_));
 sky130_fd_sc_hd__nor2_1 _2480_ (.A(_0787_),
    .B(_0813_),
    .Y(_0140_));
 sky130_fd_sc_hd__o21ai_1 _2481_ (.A1(_1245_),
    .A2(_0140_),
    .B1(_0873_),
    .Y(_0141_));
 sky130_fd_sc_hd__o311a_1 _2482_ (.A1(_0957_),
    .A2(_0767_),
    .A3(_0890_),
    .B1(_0141_),
    .C1(_0778_),
    .X(_0142_));
 sky130_fd_sc_hd__o21ba_1 _2483_ (.A1(_1356_),
    .A2(_0139_),
    .B1_N(_0142_),
    .X(_0143_));
 sky130_fd_sc_hd__a211o_1 _2484_ (.A1(_1367_),
    .A2(_0886_),
    .B1(_1112_),
    .C1(_1040_),
    .X(_0144_));
 sky130_fd_sc_hd__a311o_1 _2485_ (.A1(_1311_),
    .A2(_1219_),
    .A3(_0947_),
    .B1(_1166_),
    .C1(_1180_),
    .X(_0145_));
 sky130_fd_sc_hd__and3_2 _2486_ (.A(_0881_),
    .B(_0939_),
    .C(_0797_),
    .X(_0146_));
 sky130_fd_sc_hd__a221o_1 _2487_ (.A1(_1124_),
    .A2(_1136_),
    .B1(_1078_),
    .B2(_0806_),
    .C1(_1028_),
    .X(_0147_));
 sky130_fd_sc_hd__o311a_1 _2488_ (.A1(_1056_),
    .A2(_0980_),
    .A3(_0146_),
    .B1(_0147_),
    .C1(_0963_),
    .X(_0148_));
 sky130_fd_sc_hd__a311o_1 _2489_ (.A1(_0779_),
    .A2(_0144_),
    .A3(_0145_),
    .B1(_0148_),
    .C1(_0667_),
    .X(_0149_));
 sky130_fd_sc_hd__o21ai_4 _2490_ (.A1(_1243_),
    .A2(_0143_),
    .B1(_0149_),
    .Y(_0150_));
 sky130_fd_sc_hd__xnor2_1 _2491_ (.A(_0136_),
    .B(_0150_),
    .Y(_0151_));
 sky130_fd_sc_hd__a311o_1 _2492_ (.A1(_1367_),
    .A2(_1113_),
    .A3(_0917_),
    .B1(_1467_),
    .C1(_0725_),
    .X(_0152_));
 sky130_fd_sc_hd__or4_1 _2493_ (.A(_1060_),
    .B(_1050_),
    .C(_1190_),
    .D(_1410_),
    .X(_0153_));
 sky130_fd_sc_hd__and3_4 _2494_ (.A(_0756_),
    .B(_0745_),
    .C(_0719_),
    .X(_0154_));
 sky130_fd_sc_hd__a211o_1 _2495_ (.A1(_0806_),
    .A2(_1399_),
    .B1(_0154_),
    .C1(_0956_),
    .X(_0155_));
 sky130_fd_sc_hd__o311a_1 _2496_ (.A1(_1235_),
    .A2(_1066_),
    .A3(_1166_),
    .B1(_0155_),
    .C1(_0950_),
    .X(_0156_));
 sky130_fd_sc_hd__a31o_1 _2497_ (.A1(_1198_),
    .A2(_0152_),
    .A3(_0153_),
    .B1(_0156_),
    .X(_0157_));
 sky130_fd_sc_hd__a31o_1 _2498_ (.A1(_0852_),
    .A2(_1011_),
    .A3(_1025_),
    .B1(_0985_),
    .X(_0158_));
 sky130_fd_sc_hd__or3_1 _2499_ (.A(_0810_),
    .B(_1050_),
    .C(_1077_),
    .X(_0159_));
 sky130_fd_sc_hd__a221o_1 _2500_ (.A1(_0975_),
    .A2(_0788_),
    .B1(_1059_),
    .B2(_0881_),
    .C1(_0910_),
    .X(_0160_));
 sky130_fd_sc_hd__o311a_1 _2501_ (.A1(_1063_),
    .A2(_0733_),
    .A3(_0105_),
    .B1(_0160_),
    .C1(_0950_),
    .X(_0161_));
 sky130_fd_sc_hd__a31o_1 _2502_ (.A1(_1178_),
    .A2(_0158_),
    .A3(_0159_),
    .B1(_0161_),
    .X(_0162_));
 sky130_fd_sc_hd__and3_1 _2503_ (.A(_1041_),
    .B(_1013_),
    .C(_0738_),
    .X(_0163_));
 sky130_fd_sc_hd__and3_1 _2504_ (.A(_1117_),
    .B(_0976_),
    .C(_1073_),
    .X(_0164_));
 sky130_fd_sc_hd__or4_1 _2505_ (.A(_0984_),
    .B(_0999_),
    .C(_0814_),
    .D(_1491_),
    .X(_0165_));
 sky130_fd_sc_hd__o31a_1 _2506_ (.A1(_0725_),
    .A2(_0163_),
    .A3(_0164_),
    .B1(_0165_),
    .X(_0166_));
 sky130_fd_sc_hd__a21oi_1 _2507_ (.A1(_1113_),
    .A2(_0744_),
    .B1(_0948_),
    .Y(_0167_));
 sky130_fd_sc_hd__o221a_1 _2508_ (.A1(_0931_),
    .A2(_1008_),
    .B1(_0167_),
    .B2(_0875_),
    .C1(_0914_),
    .X(_0168_));
 sky130_fd_sc_hd__o21ba_1 _2509_ (.A1(_1198_),
    .A2(_0166_),
    .B1_N(_0168_),
    .X(_0169_));
 sky130_fd_sc_hd__or3_1 _2510_ (.A(_0810_),
    .B(_0940_),
    .C(_1084_),
    .X(_0170_));
 sky130_fd_sc_hd__or3_4 _2511_ (.A(_0836_),
    .B(_1315_),
    .C(_1277_),
    .X(_0171_));
 sky130_fd_sc_hd__nand2_2 _2512_ (.A(_1089_),
    .B(_0790_),
    .Y(_0172_));
 sky130_fd_sc_hd__and3_1 _2513_ (.A(_0716_),
    .B(_0823_),
    .C(_0790_),
    .X(_0173_));
 sky130_fd_sc_hd__a211o_1 _2514_ (.A1(_1136_),
    .A2(_0172_),
    .B1(_0173_),
    .C1(_0956_),
    .X(_0174_));
 sky130_fd_sc_hd__o311a_1 _2515_ (.A1(_1235_),
    .A2(_1127_),
    .A3(_1162_),
    .B1(_0174_),
    .C1(_0950_),
    .X(_0175_));
 sky130_fd_sc_hd__a31o_1 _2516_ (.A1(_1198_),
    .A2(_0170_),
    .A3(_0171_),
    .B1(_0175_),
    .X(_0176_));
 sky130_fd_sc_hd__mux4_2 _2517_ (.A0(_0157_),
    .A1(_0162_),
    .A2(_0169_),
    .A3(_0176_),
    .S0(_0843_),
    .S1(_0645_),
    .X(_0177_));
 sky130_fd_sc_hd__nand2_1 _2518_ (.A(_1197_),
    .B(_0177_),
    .Y(_0178_));
 sky130_fd_sc_hd__o211a_1 _2519_ (.A1(_1158_),
    .A2(_0151_),
    .B1(_0178_),
    .C1(_1242_),
    .X(_0006_));
 sky130_fd_sc_hd__a221o_1 _2520_ (.A1(_1343_),
    .A2(_0819_),
    .B1(_0976_),
    .B2(_0811_),
    .C1(_0737_),
    .X(_0179_));
 sky130_fd_sc_hd__nand2_2 _2521_ (.A(_1089_),
    .B(_0867_),
    .Y(_0180_));
 sky130_fd_sc_hd__nand2_2 _2522_ (.A(_0970_),
    .B(_0180_),
    .Y(_0181_));
 sky130_fd_sc_hd__o211a_1 _2523_ (.A1(_0743_),
    .A2(_1188_),
    .B1(_0181_),
    .C1(_0810_),
    .X(_0182_));
 sky130_fd_sc_hd__nor3_1 _2524_ (.A(_1056_),
    .B(_0893_),
    .C(_1456_),
    .Y(_0183_));
 sky130_fd_sc_hd__or3_1 _2525_ (.A(_1047_),
    .B(_0182_),
    .C(_0183_),
    .X(_0184_));
 sky130_fd_sc_hd__o211a_1 _2526_ (.A1(_1250_),
    .A2(_0179_),
    .B1(_0184_),
    .C1(_1273_),
    .X(_0185_));
 sky130_fd_sc_hd__or3_4 _2527_ (.A(_0877_),
    .B(_0887_),
    .C(_0896_),
    .X(_0186_));
 sky130_fd_sc_hd__and3_1 _2528_ (.A(_1345_),
    .B(_1344_),
    .C(_0186_),
    .X(_0187_));
 sky130_fd_sc_hd__a31o_1 _2529_ (.A1(_1403_),
    .A2(_0919_),
    .A3(_1098_),
    .B1(_1278_),
    .X(_0188_));
 sky130_fd_sc_hd__a211o_1 _2530_ (.A1(_1199_),
    .A2(net52),
    .B1(_0164_),
    .C1(_1211_),
    .X(_0189_));
 sky130_fd_sc_hd__or3_1 _2531_ (.A(_1083_),
    .B(_0827_),
    .C(_0154_),
    .X(_0190_));
 sky130_fd_sc_hd__a31o_1 _2532_ (.A1(_0703_),
    .A2(_0189_),
    .A3(_0190_),
    .B1(_1193_),
    .X(_0191_));
 sky130_fd_sc_hd__o21ba_1 _2533_ (.A1(_0187_),
    .A2(_0188_),
    .B1_N(_0191_),
    .X(_0192_));
 sky130_fd_sc_hd__or3_1 _2534_ (.A(_0645_),
    .B(_1050_),
    .C(_0146_),
    .X(_0193_));
 sky130_fd_sc_hd__o31a_1 _2535_ (.A1(_0861_),
    .A2(_0185_),
    .A3(_0192_),
    .B1(_0193_),
    .X(_0194_));
 sky130_fd_sc_hd__nor2_1 _2536_ (.A(_0771_),
    .B(_0983_),
    .Y(_0195_));
 sky130_fd_sc_hd__or3_1 _2537_ (.A(_1211_),
    .B(_0195_),
    .C(_1407_),
    .X(_0196_));
 sky130_fd_sc_hd__o311a_1 _2538_ (.A1(_1348_),
    .A2(_0720_),
    .A3(_1249_),
    .B1(_0196_),
    .C1(_1287_),
    .X(_0197_));
 sky130_fd_sc_hd__nand2_1 _2539_ (.A(_1348_),
    .B(_1174_),
    .Y(_0198_));
 sky130_fd_sc_hd__o311a_1 _2540_ (.A1(_1348_),
    .A2(_1129_),
    .A3(_0124_),
    .B1(_0198_),
    .C1(_1285_),
    .X(_0199_));
 sky130_fd_sc_hd__or2b_1 _2541_ (.A(_0762_),
    .B_N(_1107_),
    .X(_0200_));
 sky130_fd_sc_hd__a211o_2 _2542_ (.A1(_1219_),
    .A2(_1004_),
    .B1(_0890_),
    .C1(_0751_),
    .X(_0201_));
 sky130_fd_sc_hd__o21a_1 _2543_ (.A1(_0962_),
    .A2(_1530_),
    .B1(_1140_),
    .X(_0202_));
 sky130_fd_sc_hd__o211a_1 _2544_ (.A1(_0737_),
    .A2(_1011_),
    .B1(_0093_),
    .C1(_0922_),
    .X(_0203_));
 sky130_fd_sc_hd__o21a_2 _2545_ (.A1(_0202_),
    .A2(_0203_),
    .B1(_1115_),
    .X(_0204_));
 sky130_fd_sc_hd__a311o_1 _2546_ (.A1(_0779_),
    .A2(_0200_),
    .A3(_0201_),
    .B1(_0204_),
    .C1(_0667_),
    .X(_0205_));
 sky130_fd_sc_hd__o311a_1 _2547_ (.A1(_1273_),
    .A2(_0197_),
    .A3(_0199_),
    .B1(_0205_),
    .C1(_1396_),
    .X(_0206_));
 sky130_fd_sc_hd__or4_1 _2548_ (.A(_1049_),
    .B(_0733_),
    .C(_1183_),
    .D(_1265_),
    .X(_0207_));
 sky130_fd_sc_hd__o311a_1 _2549_ (.A1(_1348_),
    .A2(_0733_),
    .A3(_1524_),
    .B1(_0207_),
    .C1(_1310_),
    .X(_0208_));
 sky130_fd_sc_hd__and2_2 _2550_ (.A(_0758_),
    .B(_0976_),
    .X(_0209_));
 sky130_fd_sc_hd__a221o_1 _2551_ (.A1(_1367_),
    .A2(_0886_),
    .B1(_0961_),
    .B2(_0829_),
    .C1(_1264_),
    .X(_0210_));
 sky130_fd_sc_hd__o311a_1 _2552_ (.A1(_1403_),
    .A2(_1300_),
    .A3(_0209_),
    .B1(_0210_),
    .C1(_1356_),
    .X(_0211_));
 sky130_fd_sc_hd__or3_1 _2553_ (.A(_0936_),
    .B(_1077_),
    .C(_0137_),
    .X(_0212_));
 sky130_fd_sc_hd__or3_1 _2554_ (.A(_0725_),
    .B(_0938_),
    .C(_0154_),
    .X(_0213_));
 sky130_fd_sc_hd__and2_1 _2555_ (.A(_1106_),
    .B(_1254_),
    .X(_0214_));
 sky130_fd_sc_hd__or3b_4 _2556_ (.A(_0724_),
    .B(_0832_),
    .C_N(_1214_),
    .X(_0215_));
 sky130_fd_sc_hd__o311a_1 _2557_ (.A1(_0945_),
    .A2(_1175_),
    .A3(_0214_),
    .B1(_0215_),
    .C1(_0978_),
    .X(_0216_));
 sky130_fd_sc_hd__a311o_1 _2558_ (.A1(_1310_),
    .A2(_0212_),
    .A3(_0213_),
    .B1(_0216_),
    .C1(_1318_),
    .X(_0217_));
 sky130_fd_sc_hd__o311a_1 _2559_ (.A1(_1298_),
    .A2(_0208_),
    .A3(_0211_),
    .B1(_0217_),
    .C1(_0861_),
    .X(_0218_));
 sky130_fd_sc_hd__o21ai_1 _2560_ (.A1(_0206_),
    .A2(_0218_),
    .B1(_1197_),
    .Y(_0219_));
 sky130_fd_sc_hd__o211a_1 _2561_ (.A1(_1158_),
    .A2(_0194_),
    .B1(_0219_),
    .C1(_1242_),
    .X(_0007_));
 sky130_fd_sc_hd__and3_1 _2562_ (.A(_0860_),
    .B(_0803_),
    .C(_1020_),
    .X(_0220_));
 sky130_fd_sc_hd__and3_2 _2563_ (.A(_0770_),
    .B(_1019_),
    .C(_0983_),
    .X(_0221_));
 sky130_fd_sc_hd__a221o_1 _2564_ (.A1(_0824_),
    .A2(_0827_),
    .B1(_1099_),
    .B2(_0803_),
    .C1(_1235_),
    .X(_0222_));
 sky130_fd_sc_hd__o311a_1 _2565_ (.A1(_0811_),
    .A2(_1470_),
    .A3(_0221_),
    .B1(_0222_),
    .C1(_0907_),
    .X(_0223_));
 sky130_fd_sc_hd__or3_1 _2566_ (.A(_0755_),
    .B(_0966_),
    .C(_1305_),
    .X(_0224_));
 sky130_fd_sc_hd__o311a_1 _2567_ (.A1(_1256_),
    .A2(_0931_),
    .A3(_0146_),
    .B1(_0224_),
    .C1(_1193_),
    .X(_0225_));
 sky130_fd_sc_hd__a211o_1 _2568_ (.A1(_0824_),
    .A2(_0815_),
    .B1(_1475_),
    .C1(_1211_),
    .X(_0226_));
 sky130_fd_sc_hd__a21o_1 _2569_ (.A1(_0917_),
    .A2(_1066_),
    .B1(_0942_),
    .X(_0227_));
 sky130_fd_sc_hd__or3b_1 _2570_ (.A(_0864_),
    .B(_1026_),
    .C_N(_1065_),
    .X(_0228_));
 sky130_fd_sc_hd__o311a_1 _2571_ (.A1(_1063_),
    .A2(_1141_),
    .A3(_1302_),
    .B1(_0228_),
    .C1(_0661_),
    .X(_0229_));
 sky130_fd_sc_hd__a311o_1 _2572_ (.A1(_1193_),
    .A2(_0226_),
    .A3(_0227_),
    .B1(_1178_),
    .C1(_0229_),
    .X(_0230_));
 sky130_fd_sc_hd__o31a_2 _2573_ (.A1(_0706_),
    .A2(_0223_),
    .A3(_0225_),
    .B1(_0230_),
    .X(_0231_));
 sky130_fd_sc_hd__xnor2_1 _2574_ (.A(_0220_),
    .B(_0231_),
    .Y(_0232_));
 sky130_fd_sc_hd__or3_1 _2575_ (.A(_0936_),
    .B(_1162_),
    .C(_1288_),
    .X(_0233_));
 sky130_fd_sc_hd__o311a_1 _2576_ (.A1(_1403_),
    .A2(_1174_),
    .A3(_1432_),
    .B1(_0233_),
    .C1(_1308_),
    .X(_0234_));
 sky130_fd_sc_hd__o221a_1 _2577_ (.A1(_1259_),
    .A2(_1004_),
    .B1(_1112_),
    .B2(_1151_),
    .C1(_1285_),
    .X(_0235_));
 sky130_fd_sc_hd__a311o_1 _2578_ (.A1(_1089_),
    .A2(_1199_),
    .A3(_1019_),
    .B1(_1276_),
    .C1(_1109_),
    .X(_0236_));
 sky130_fd_sc_hd__nor2_1 _2579_ (.A(_0760_),
    .B(_0867_),
    .Y(_0237_));
 sky130_fd_sc_hd__o21ai_1 _2580_ (.A1(_0237_),
    .A2(_1379_),
    .B1(_1335_),
    .Y(_0238_));
 sky130_fd_sc_hd__a211o_1 _2581_ (.A1(_0803_),
    .A2(_1072_),
    .B1(_0146_),
    .C1(_0985_),
    .X(_0239_));
 sky130_fd_sc_hd__o311a_1 _2582_ (.A1(_0957_),
    .A2(_1326_),
    .A3(_1501_),
    .B1(_0239_),
    .C1(_0778_),
    .X(_0240_));
 sky130_fd_sc_hd__a311o_1 _2583_ (.A1(_1310_),
    .A2(_0236_),
    .A3(_0238_),
    .B1(_0240_),
    .C1(_1318_),
    .X(_0241_));
 sky130_fd_sc_hd__o31ai_2 _2584_ (.A1(_1298_),
    .A2(_0234_),
    .A3(_0235_),
    .B1(_0241_),
    .Y(_0242_));
 sky130_fd_sc_hd__a221o_1 _2585_ (.A1(_1013_),
    .A2(_1206_),
    .B1(_0180_),
    .B2(_1011_),
    .C1(_0800_),
    .X(_0243_));
 sky130_fd_sc_hd__o311a_1 _2586_ (.A1(_1109_),
    .A2(_0925_),
    .A3(_1354_),
    .B1(_0243_),
    .C1(_0978_),
    .X(_0244_));
 sky130_fd_sc_hd__a311o_1 _2587_ (.A1(_0878_),
    .A2(_0713_),
    .A3(_0971_),
    .B1(_1166_),
    .C1(_1060_),
    .X(_0245_));
 sky130_fd_sc_hd__o311a_1 _2588_ (.A1(_0751_),
    .A2(_1294_),
    .A3(_1500_),
    .B1(_0245_),
    .C1(_1047_),
    .X(_0246_));
 sky130_fd_sc_hd__or3_1 _2589_ (.A(_0800_),
    .B(_1119_),
    .C(_1467_),
    .X(_0247_));
 sky130_fd_sc_hd__o311a_1 _2590_ (.A1(_1165_),
    .A2(_1229_),
    .A3(_1072_),
    .B1(_0247_),
    .C1(_0839_),
    .X(_0248_));
 sky130_fd_sc_hd__a22o_1 _2591_ (.A1(_0769_),
    .A2(_0989_),
    .B1(_1325_),
    .B2(_0854_),
    .X(_0249_));
 sky130_fd_sc_hd__a21o_1 _2592_ (.A1(_1065_),
    .A2(_0249_),
    .B1(_1063_),
    .X(_0250_));
 sky130_fd_sc_hd__a211o_1 _2593_ (.A1(_1000_),
    .A2(_0815_),
    .B1(_1266_),
    .C1(_1049_),
    .X(_0251_));
 sky130_fd_sc_hd__a31o_1 _2594_ (.A1(_0915_),
    .A2(_0250_),
    .A3(_0251_),
    .B1(_0842_),
    .X(_0252_));
 sky130_fd_sc_hd__o32a_2 _2595_ (.A1(_0667_),
    .A2(_0244_),
    .A3(_0246_),
    .B1(_0248_),
    .B2(_0252_),
    .X(_0253_));
 sky130_fd_sc_hd__nor2_1 _2596_ (.A(_0861_),
    .B(_0253_),
    .Y(_0254_));
 sky130_fd_sc_hd__a211o_1 _2597_ (.A1(_1365_),
    .A2(_0242_),
    .B1(_0254_),
    .C1(_1322_),
    .X(_0255_));
 sky130_fd_sc_hd__o211a_1 _2598_ (.A1(_1158_),
    .A2(_0232_),
    .B1(_0255_),
    .C1(_1242_),
    .X(_0008_));
 sky130_fd_sc_hd__nand2_1 _2599_ (.A(_0878_),
    .B(_0989_),
    .Y(_0256_));
 sky130_fd_sc_hd__or3_2 _2600_ (.A(_0715_),
    .B(_0998_),
    .C(_0818_),
    .X(_0257_));
 sky130_fd_sc_hd__nor2_1 _2601_ (.A(_0751_),
    .B(_0928_),
    .Y(_0258_));
 sky130_fd_sc_hd__a32o_1 _2602_ (.A1(_0811_),
    .A2(_1160_),
    .A3(_0256_),
    .B1(_0257_),
    .B2(_0258_),
    .X(_0259_));
 sky130_fd_sc_hd__o221a_1 _2603_ (.A1(_0869_),
    .A2(_1236_),
    .B1(_1399_),
    .B2(_0770_),
    .C1(_0810_),
    .X(_0260_));
 sky130_fd_sc_hd__a311o_1 _2604_ (.A1(_1256_),
    .A2(_1214_),
    .A3(_0257_),
    .B1(_0260_),
    .C1(_0915_),
    .X(_0261_));
 sky130_fd_sc_hd__o211a_1 _2605_ (.A1(_1342_),
    .A2(_0259_),
    .B1(_0261_),
    .C1(_0843_),
    .X(_0262_));
 sky130_fd_sc_hd__o221a_1 _2606_ (.A1(_1343_),
    .A2(_0195_),
    .B1(_1001_),
    .B2(_1124_),
    .C1(_1291_),
    .X(_0263_));
 sky130_fd_sc_hd__nand2_1 _2607_ (.A(_1206_),
    .B(_1025_),
    .Y(_0264_));
 sky130_fd_sc_hd__a31o_1 _2608_ (.A1(_1256_),
    .A2(_1453_),
    .A3(_0264_),
    .B1(_0839_),
    .X(_0265_));
 sky130_fd_sc_hd__and3_2 _2609_ (.A(_0939_),
    .B(_0738_),
    .C(_0924_),
    .X(_0266_));
 sky130_fd_sc_hd__o21ai_1 _2610_ (.A1(_1030_),
    .A2(_0266_),
    .B1(_1165_),
    .Y(_0267_));
 sky130_fd_sc_hd__o31a_1 _2611_ (.A1(_1165_),
    .A2(_1206_),
    .A3(_1466_),
    .B1(_0267_),
    .X(_0268_));
 sky130_fd_sc_hd__o221a_1 _2612_ (.A1(_0263_),
    .A2(_0265_),
    .B1(_0268_),
    .B2(_1250_),
    .C1(_1164_),
    .X(_0269_));
 sky130_fd_sc_hd__and3_1 _2613_ (.A(_0770_),
    .B(_1219_),
    .C(_0976_),
    .X(_0270_));
 sky130_fd_sc_hd__o21ai_1 _2614_ (.A1(_1366_),
    .A2(_0270_),
    .B1(_1345_),
    .Y(_0271_));
 sky130_fd_sc_hd__o31a_1 _2615_ (.A1(_1281_),
    .A2(_0974_),
    .A3(_1443_),
    .B1(_0271_),
    .X(_0272_));
 sky130_fd_sc_hd__nor2_2 _2616_ (.A(_1136_),
    .B(_1213_),
    .Y(_0273_));
 sky130_fd_sc_hd__a311o_1 _2617_ (.A1(_1232_),
    .A2(_0786_),
    .A3(_0867_),
    .B1(_0273_),
    .C1(_0873_),
    .X(_0274_));
 sky130_fd_sc_hd__or4_1 _2618_ (.A(_1060_),
    .B(_1030_),
    .C(_0997_),
    .D(_1314_),
    .X(_0275_));
 sky130_fd_sc_hd__a31o_1 _2619_ (.A1(_1198_),
    .A2(_0274_),
    .A3(_0275_),
    .B1(_0907_),
    .X(_0276_));
 sky130_fd_sc_hd__o21ba_1 _2620_ (.A1(_1250_),
    .A2(_0272_),
    .B1_N(_0276_),
    .X(_0277_));
 sky130_fd_sc_hd__o21ai_1 _2621_ (.A1(_1199_),
    .A2(_1506_),
    .B1(_0080_),
    .Y(_0278_));
 sky130_fd_sc_hd__and3_1 _2622_ (.A(_0873_),
    .B(_0854_),
    .C(_0739_),
    .X(_0279_));
 sky130_fd_sc_hd__nor2_1 _2623_ (.A(_1261_),
    .B(_0278_),
    .Y(_0280_));
 sky130_fd_sc_hd__a211o_2 _2624_ (.A1(_0278_),
    .A2(_0279_),
    .B1(_0280_),
    .C1(_1278_),
    .X(_0281_));
 sky130_fd_sc_hd__and3b_1 _2625_ (.A_N(_1255_),
    .B(_1049_),
    .C(_0722_),
    .X(_0282_));
 sky130_fd_sc_hd__a221o_1 _2626_ (.A1(_0786_),
    .A2(_0965_),
    .B1(_1399_),
    .B2(_0807_),
    .C1(_0836_),
    .X(_0283_));
 sky130_fd_sc_hd__or3b_1 _2627_ (.A(_0915_),
    .B(_0282_),
    .C_N(_0283_),
    .X(_0284_));
 sky130_fd_sc_hd__a31o_1 _2628_ (.A1(_1164_),
    .A2(_0281_),
    .A3(_0284_),
    .B1(_1039_),
    .X(_0285_));
 sky130_fd_sc_hd__o32a_1 _2629_ (.A1(_1396_),
    .A2(_0262_),
    .A3(_0269_),
    .B1(_0277_),
    .B2(_0285_),
    .X(_0286_));
 sky130_fd_sc_hd__o21ai_1 _2630_ (.A1(_0983_),
    .A2(_1314_),
    .B1(_1335_),
    .Y(_0287_));
 sky130_fd_sc_hd__o311a_1 _2631_ (.A1(_1345_),
    .A2(_0798_),
    .A3(_1512_),
    .B1(_0287_),
    .C1(_0935_),
    .X(_0288_));
 sky130_fd_sc_hd__and3_1 _2632_ (.A(_0820_),
    .B(_0924_),
    .C(_0947_),
    .X(_0289_));
 sky130_fd_sc_hd__a21o_1 _2633_ (.A1(_1347_),
    .A2(_1097_),
    .B1(_1259_),
    .X(_0290_));
 sky130_fd_sc_hd__o311a_1 _2634_ (.A1(_1348_),
    .A2(_1079_),
    .A3(_0289_),
    .B1(_0290_),
    .C1(_1310_),
    .X(_0291_));
 sky130_fd_sc_hd__a22o_1 _2635_ (.A1(_0970_),
    .A2(_1506_),
    .B1(_1324_),
    .B2(_0929_),
    .X(_0292_));
 sky130_fd_sc_hd__nor2_1 _2636_ (.A(_1247_),
    .B(_0289_),
    .Y(_0293_));
 sky130_fd_sc_hd__mux2_1 _2637_ (.A0(_0292_),
    .A1(_0293_),
    .S(_0957_),
    .X(_0294_));
 sky130_fd_sc_hd__a211o_1 _2638_ (.A1(_0878_),
    .A2(_0973_),
    .B1(_0130_),
    .C1(_0922_),
    .X(_0295_));
 sky130_fd_sc_hd__o311a_1 _2639_ (.A1(_1109_),
    .A2(_1236_),
    .A3(_1523_),
    .B1(_0295_),
    .C1(_0782_),
    .X(_0296_));
 sky130_fd_sc_hd__a211o_1 _2640_ (.A1(_1342_),
    .A2(_0294_),
    .B1(_0296_),
    .C1(_0952_),
    .X(_0297_));
 sky130_fd_sc_hd__o311a_2 _2641_ (.A1(_0673_),
    .A2(_0288_),
    .A3(_0291_),
    .B1(_0297_),
    .C1(_1161_),
    .X(_0298_));
 sky130_fd_sc_hd__a21oi_1 _2642_ (.A1(_0871_),
    .A2(_1065_),
    .B1(_0655_),
    .Y(_0299_));
 sky130_fd_sc_hd__o21ai_1 _2643_ (.A1(_0298_),
    .A2(_0299_),
    .B1(_1322_),
    .Y(_0300_));
 sky130_fd_sc_hd__o211a_1 _2644_ (.A1(_1322_),
    .A2(_0286_),
    .B1(_0300_),
    .C1(_1242_),
    .X(_0009_));
 sky130_fd_sc_hd__a211o_1 _2645_ (.A1(_1124_),
    .A2(_0816_),
    .B1(_1142_),
    .C1(_1281_),
    .X(_0301_));
 sky130_fd_sc_hd__or3_1 _2646_ (.A(_0811_),
    .B(_0154_),
    .C(_0173_),
    .X(_0302_));
 sky130_fd_sc_hd__and3_2 _2647_ (.A(_0741_),
    .B(_0728_),
    .C(net54),
    .X(_0303_));
 sky130_fd_sc_hd__or3_1 _2648_ (.A(_1235_),
    .B(_1380_),
    .C(_1511_),
    .X(_0304_));
 sky130_fd_sc_hd__o211a_1 _2649_ (.A1(_1147_),
    .A2(_0303_),
    .B1(_0304_),
    .C1(_0935_),
    .X(_0305_));
 sky130_fd_sc_hd__a311o_1 _2650_ (.A1(_0706_),
    .A2(_0301_),
    .A3(_0302_),
    .B1(_0305_),
    .C1(_1164_),
    .X(_0306_));
 sky130_fd_sc_hd__or3_1 _2651_ (.A(_1083_),
    .B(_1009_),
    .C(_0266_),
    .X(_0307_));
 sky130_fd_sc_hd__o311a_1 _2652_ (.A1(_1256_),
    .A2(_1475_),
    .A3(net52),
    .B1(_0307_),
    .C1(_0703_),
    .X(_0308_));
 sky130_fd_sc_hd__nor2_1 _2653_ (.A(_1016_),
    .B(_1301_),
    .Y(_0309_));
 sky130_fd_sc_hd__o221a_1 _2654_ (.A1(_0816_),
    .A2(_1500_),
    .B1(_0309_),
    .B2(_1274_),
    .C1(_1178_),
    .X(_0310_));
 sky130_fd_sc_hd__or3_1 _2655_ (.A(_0843_),
    .B(_0308_),
    .C(_0310_),
    .X(_0311_));
 sky130_fd_sc_hd__a21oi_1 _2656_ (.A1(_0306_),
    .A2(_0311_),
    .B1(_1365_),
    .Y(_0312_));
 sky130_fd_sc_hd__nor2_1 _2657_ (.A(_0655_),
    .B(_0989_),
    .Y(_0313_));
 sky130_fd_sc_hd__o31ai_1 _2658_ (.A1(_0720_),
    .A2(_0901_),
    .A3(_1314_),
    .B1(_1256_),
    .Y(_0314_));
 sky130_fd_sc_hd__o311a_1 _2659_ (.A1(_1345_),
    .A2(_1129_),
    .A3(_0209_),
    .B1(_0314_),
    .C1(_1287_),
    .X(_0315_));
 sky130_fd_sc_hd__nand2_1 _2660_ (.A(_1261_),
    .B(_1329_),
    .Y(_0316_));
 sky130_fd_sc_hd__a211o_1 _2661_ (.A1(_1073_),
    .A2(_1379_),
    .B1(_1137_),
    .C1(_0801_),
    .X(_0317_));
 sky130_fd_sc_hd__o211a_1 _2662_ (.A1(_0977_),
    .A2(_0316_),
    .B1(_0317_),
    .C1(_1285_),
    .X(_0318_));
 sky130_fd_sc_hd__or4_1 _2663_ (.A(_0755_),
    .B(_0805_),
    .C(_1016_),
    .D(_1330_),
    .X(_0319_));
 sky130_fd_sc_hd__o21ai_1 _2664_ (.A1(_1190_),
    .A2(_1456_),
    .B1(_1274_),
    .Y(_0320_));
 sky130_fd_sc_hd__or3_1 _2665_ (.A(_0835_),
    .B(_0733_),
    .C(_0855_),
    .X(_0321_));
 sky130_fd_sc_hd__o311a_1 _2666_ (.A1(_1056_),
    .A2(_0903_),
    .A3(_1379_),
    .B1(_0321_),
    .C1(_0778_),
    .X(_0322_));
 sky130_fd_sc_hd__a311o_1 _2667_ (.A1(_1287_),
    .A2(_0319_),
    .A3(_0320_),
    .B1(_0322_),
    .C1(_0667_),
    .X(_0323_));
 sky130_fd_sc_hd__o311a_1 _2668_ (.A1(_1273_),
    .A2(_0315_),
    .A3(_0318_),
    .B1(_0323_),
    .C1(_1161_),
    .X(_0324_));
 sky130_fd_sc_hd__a221o_1 _2669_ (.A1(_1000_),
    .A2(_0917_),
    .B1(_0819_),
    .B2(_1311_),
    .C1(_1180_),
    .X(_0325_));
 sky130_fd_sc_hd__o311a_1 _2670_ (.A1(_1345_),
    .A2(_0960_),
    .A3(_1059_),
    .B1(_0325_),
    .C1(_1287_),
    .X(_0326_));
 sky130_fd_sc_hd__a221o_1 _2671_ (.A1(_1311_),
    .A2(_1097_),
    .B1(_1127_),
    .B2(_0824_),
    .C1(_1264_),
    .X(_0327_));
 sky130_fd_sc_hd__o311a_1 _2672_ (.A1(_1403_),
    .A2(_1088_),
    .A3(_1027_),
    .B1(_0327_),
    .C1(_1285_),
    .X(_0328_));
 sky130_fd_sc_hd__or3b_1 _2673_ (.A(_0873_),
    .B(_0747_),
    .C_N(_1065_),
    .X(_0329_));
 sky130_fd_sc_hd__nand3_1 _2674_ (.A(_1274_),
    .B(_0871_),
    .C(_0181_),
    .Y(_0330_));
 sky130_fd_sc_hd__and3_1 _2675_ (.A(_0926_),
    .B(_0713_),
    .C(_0892_),
    .X(_0331_));
 sky130_fd_sc_hd__a311o_1 _2676_ (.A1(_1136_),
    .A2(_0854_),
    .A3(_1325_),
    .B1(_0331_),
    .C1(_0750_),
    .X(_0332_));
 sky130_fd_sc_hd__o311a_1 _2677_ (.A1(_0945_),
    .A2(_0747_),
    .A3(_1027_),
    .B1(_0332_),
    .C1(_0778_),
    .X(_0333_));
 sky130_fd_sc_hd__a311o_1 _2678_ (.A1(_1287_),
    .A2(_0329_),
    .A3(_0330_),
    .B1(_0333_),
    .C1(_1318_),
    .X(_0334_));
 sky130_fd_sc_hd__o311a_1 _2679_ (.A1(_1298_),
    .A2(_0326_),
    .A3(_0328_),
    .B1(_0334_),
    .C1(_1039_),
    .X(_0335_));
 sky130_fd_sc_hd__o21ai_1 _2680_ (.A1(_0324_),
    .A2(_0335_),
    .B1(_1197_),
    .Y(_0336_));
 sky130_fd_sc_hd__o311a_1 _2681_ (.A1(_1158_),
    .A2(_0312_),
    .A3(_0313_),
    .B1(_0336_),
    .C1(_0859_),
    .X(_0010_));
 sky130_fd_sc_hd__and2b_1 _2682_ (.A_N(_0900_),
    .B(_1003_),
    .X(_0337_));
 sky130_fd_sc_hd__o311a_1 _2683_ (.A1(_0771_),
    .A2(_1347_),
    .A3(_0760_),
    .B1(_1453_),
    .C1(_1274_),
    .X(_0338_));
 sky130_fd_sc_hd__a21oi_1 _2684_ (.A1(_1067_),
    .A2(_1519_),
    .B1(_1291_),
    .Y(_0339_));
 sky130_fd_sc_hd__nor2_4 _2685_ (.A(_0756_),
    .B(_0760_),
    .Y(_0340_));
 sky130_fd_sc_hd__o221a_1 _2686_ (.A1(_0852_),
    .A2(_1311_),
    .B1(_0340_),
    .B2(_1300_),
    .C1(_0923_),
    .X(_0341_));
 sky130_fd_sc_hd__o21ai_1 _2687_ (.A1(_0339_),
    .A2(_0341_),
    .B1(_0783_),
    .Y(_0342_));
 sky130_fd_sc_hd__o31a_1 _2688_ (.A1(_0783_),
    .A2(_0337_),
    .A3(_0338_),
    .B1(_0342_),
    .X(_0343_));
 sky130_fd_sc_hd__and3_1 _2689_ (.A(_1232_),
    .B(_1041_),
    .C(_1025_),
    .X(_0344_));
 sky130_fd_sc_hd__and3_2 _2690_ (.A(_0939_),
    .B(_0831_),
    .C(_0897_),
    .X(_0345_));
 sky130_fd_sc_hd__or3_1 _2691_ (.A(_0873_),
    .B(_0344_),
    .C(_0345_),
    .X(_0346_));
 sky130_fd_sc_hd__o311a_1 _2692_ (.A1(_1299_),
    .A2(_1302_),
    .A3(_1417_),
    .B1(_0346_),
    .C1(_0779_),
    .X(_0347_));
 sky130_fd_sc_hd__a221o_1 _2693_ (.A1(_1000_),
    .A2(_0816_),
    .B1(_1023_),
    .B2(_1219_),
    .C1(_1264_),
    .X(_0348_));
 sky130_fd_sc_hd__o311a_1 _2694_ (.A1(_1403_),
    .A2(_0948_),
    .A3(_1002_),
    .B1(_0348_),
    .C1(_1308_),
    .X(_0349_));
 sky130_fd_sc_hd__o21ai_2 _2695_ (.A1(_0347_),
    .A2(_0349_),
    .B1(_1243_),
    .Y(_0350_));
 sky130_fd_sc_hd__o211a_1 _2696_ (.A1(_1243_),
    .A2(_0343_),
    .B1(_0350_),
    .C1(_0655_),
    .X(_0351_));
 sky130_fd_sc_hd__a211oi_1 _2697_ (.A1(_1347_),
    .A2(_1254_),
    .B1(net51),
    .C1(_0655_),
    .Y(_0352_));
 sky130_fd_sc_hd__nand2_1 _2698_ (.A(_0755_),
    .B(_1167_),
    .Y(_0353_));
 sky130_fd_sc_hd__o31a_1 _2699_ (.A1(_1180_),
    .A2(_0829_),
    .A3(_1135_),
    .B1(_0963_),
    .X(_0354_));
 sky130_fd_sc_hd__o21a_1 _2700_ (.A1(_1410_),
    .A2(_0353_),
    .B1(_0354_),
    .X(_0355_));
 sky130_fd_sc_hd__a211o_1 _2701_ (.A1(_1367_),
    .A2(_0973_),
    .B1(_1410_),
    .C1(_0801_),
    .X(_0356_));
 sky130_fd_sc_hd__o311a_1 _2702_ (.A1(_1281_),
    .A2(_1300_),
    .A3(_0214_),
    .B1(_0356_),
    .C1(_1285_),
    .X(_0357_));
 sky130_fd_sc_hd__or2_1 _2703_ (.A(_0834_),
    .B(_0899_),
    .X(_0358_));
 sky130_fd_sc_hd__a22o_1 _2704_ (.A1(_0880_),
    .A2(_1016_),
    .B1(_1073_),
    .B2(_1077_),
    .X(_0359_));
 sky130_fd_sc_hd__a2bb2o_1 _2705_ (.A1_N(_0273_),
    .A2_N(_0358_),
    .B1(_0359_),
    .B2(_1264_),
    .X(_0360_));
 sky130_fd_sc_hd__a211o_1 _2706_ (.A1(_0999_),
    .A2(_0815_),
    .B1(_1183_),
    .C1(_1028_),
    .X(_0361_));
 sky130_fd_sc_hd__a21o_1 _2707_ (.A1(_0791_),
    .A2(_1358_),
    .B1(_0922_),
    .X(_0362_));
 sky130_fd_sc_hd__and3_1 _2708_ (.A(_0963_),
    .B(_0361_),
    .C(_0362_),
    .X(_0363_));
 sky130_fd_sc_hd__a211o_1 _2709_ (.A1(_1356_),
    .A2(_0360_),
    .B1(_0363_),
    .C1(_0860_),
    .X(_0364_));
 sky130_fd_sc_hd__o311a_1 _2710_ (.A1(_0645_),
    .A2(_0355_),
    .A3(_0357_),
    .B1(_0364_),
    .C1(_0673_),
    .X(_0365_));
 sky130_fd_sc_hd__o21ai_1 _2711_ (.A1(_1125_),
    .A2(_1334_),
    .B1(_1335_),
    .Y(_0366_));
 sky130_fd_sc_hd__o311a_1 _2712_ (.A1(_0787_),
    .A2(_1259_),
    .A3(_1044_),
    .B1(_0366_),
    .C1(_0779_),
    .X(_0367_));
 sky130_fd_sc_hd__a221o_1 _2713_ (.A1(_1367_),
    .A2(_0824_),
    .B1(_0807_),
    .B2(_1020_),
    .C1(_1040_),
    .X(_0368_));
 sky130_fd_sc_hd__o311a_1 _2714_ (.A1(_1403_),
    .A2(_1079_),
    .A3(_0154_),
    .B1(_0368_),
    .C1(_1308_),
    .X(_0369_));
 sky130_fd_sc_hd__a221o_1 _2715_ (.A1(_1013_),
    .A2(_0827_),
    .B1(_0929_),
    .B2(_0960_),
    .C1(_0964_),
    .X(_0370_));
 sky130_fd_sc_hd__o311a_1 _2716_ (.A1(_0873_),
    .A2(_0805_),
    .A3(_0273_),
    .B1(_0370_),
    .C1(_0934_),
    .X(_0371_));
 sky130_fd_sc_hd__a211o_1 _2717_ (.A1(_0916_),
    .A2(_1152_),
    .B1(_0266_),
    .C1(_0750_),
    .X(_0372_));
 sky130_fd_sc_hd__o211a_1 _2718_ (.A1(_1109_),
    .A2(_0902_),
    .B1(_0372_),
    .C1(_0963_),
    .X(_0373_));
 sky130_fd_sc_hd__or3_1 _2719_ (.A(_0634_),
    .B(_0371_),
    .C(_0373_),
    .X(_0374_));
 sky130_fd_sc_hd__o311a_1 _2720_ (.A1(_1039_),
    .A2(_0367_),
    .A3(_0369_),
    .B1(_0374_),
    .C1(_1243_),
    .X(_0375_));
 sky130_fd_sc_hd__o21ai_1 _2721_ (.A1(_0365_),
    .A2(_0375_),
    .B1(_1197_),
    .Y(_0376_));
 sky130_fd_sc_hd__o311a_1 _2722_ (.A1(_1158_),
    .A2(_0351_),
    .A3(_0352_),
    .B1(_0376_),
    .C1(_0859_),
    .X(_0011_));
 sky130_fd_sc_hd__o21a_1 _2723_ (.A1(_1347_),
    .A2(_0903_),
    .B1(_0919_),
    .X(_0377_));
 sky130_fd_sc_hd__or3_1 _2724_ (.A(_0911_),
    .B(_0974_),
    .C(_1094_),
    .X(_0378_));
 sky130_fd_sc_hd__o211a_1 _2725_ (.A1(_0752_),
    .A2(_0377_),
    .B1(_0378_),
    .C1(_0783_),
    .X(_0379_));
 sky130_fd_sc_hd__nor2_2 _2726_ (.A(_0771_),
    .B(_0896_),
    .Y(_0380_));
 sky130_fd_sc_hd__o21ai_1 _2727_ (.A1(_1438_),
    .A2(_0221_),
    .B1(_1244_),
    .Y(_0381_));
 sky130_fd_sc_hd__o311a_1 _2728_ (.A1(_1244_),
    .A2(_0380_),
    .A3(_1125_),
    .B1(_0381_),
    .C1(_1342_),
    .X(_0382_));
 sky130_fd_sc_hd__o21ai_1 _2729_ (.A1(_1252_),
    .A2(_1334_),
    .B1(_0752_),
    .Y(_0383_));
 sky130_fd_sc_hd__o31a_1 _2730_ (.A1(_1391_),
    .A2(_0744_),
    .A3(_1147_),
    .B1(_0915_),
    .X(_0384_));
 sky130_fd_sc_hd__o211a_1 _2731_ (.A1(_1199_),
    .A2(_0340_),
    .B1(_0256_),
    .C1(_1211_),
    .X(_0385_));
 sky130_fd_sc_hd__a31o_1 _2732_ (.A1(_1291_),
    .A2(_0181_),
    .A3(_0186_),
    .B1(_0385_),
    .X(_0386_));
 sky130_fd_sc_hd__a221o_1 _2733_ (.A1(_0383_),
    .A2(_0384_),
    .B1(_0386_),
    .B2(_1342_),
    .C1(_0843_),
    .X(_0387_));
 sky130_fd_sc_hd__o311a_1 _2734_ (.A1(_0673_),
    .A2(_0379_),
    .A3(_0382_),
    .B1(_0387_),
    .C1(_0655_),
    .X(_0388_));
 sky130_fd_sc_hd__nor2_2 _2735_ (.A(_1123_),
    .B(_0877_),
    .Y(_0389_));
 sky130_fd_sc_hd__nand2_1 _2736_ (.A(_0806_),
    .B(_0867_),
    .Y(_0390_));
 sky130_fd_sc_hd__a21o_1 _2737_ (.A1(_0390_),
    .A2(_0983_),
    .B1(_1261_),
    .X(_0391_));
 sky130_fd_sc_hd__o311a_1 _2738_ (.A1(_1281_),
    .A2(_0807_),
    .A3(_0389_),
    .B1(_0391_),
    .C1(_1285_),
    .X(_0392_));
 sky130_fd_sc_hd__a21oi_1 _2739_ (.A1(_0452_),
    .A2(_0813_),
    .B1(_0720_),
    .Y(_0393_));
 sky130_fd_sc_hd__o221a_1 _2740_ (.A1(_1299_),
    .A2(_1323_),
    .B1(_0393_),
    .B2(_0752_),
    .C1(_1308_),
    .X(_0394_));
 sky130_fd_sc_hd__a221o_1 _2741_ (.A1(_1124_),
    .A2(_1229_),
    .B1(_1072_),
    .B2(_0803_),
    .C1(_1261_),
    .X(_0395_));
 sky130_fd_sc_hd__o311a_1 _2742_ (.A1(_1244_),
    .A2(_1072_),
    .A3(_0109_),
    .B1(_0395_),
    .C1(_0783_),
    .X(_0396_));
 sky130_fd_sc_hd__o21ai_1 _2743_ (.A1(_1190_),
    .A2(_0214_),
    .B1(_1244_),
    .Y(_0397_));
 sky130_fd_sc_hd__a21o_1 _2744_ (.A1(_1229_),
    .A2(_1399_),
    .B1(_1259_),
    .X(_0398_));
 sky130_fd_sc_hd__a31o_1 _2745_ (.A1(_1342_),
    .A2(_0397_),
    .A3(_0398_),
    .B1(_0952_),
    .X(_0399_));
 sky130_fd_sc_hd__o32a_1 _2746_ (.A1(_0673_),
    .A2(_0392_),
    .A3(_0394_),
    .B1(_0396_),
    .B2(_0399_),
    .X(_0400_));
 sky130_fd_sc_hd__nor2_1 _2747_ (.A(_0655_),
    .B(_0400_),
    .Y(_0401_));
 sky130_fd_sc_hd__nand2_1 _2748_ (.A(_0929_),
    .B(_1206_),
    .Y(_0402_));
 sky130_fd_sc_hd__a211o_1 _2749_ (.A1(_0917_),
    .A2(_1045_),
    .B1(_1189_),
    .C1(_0957_),
    .X(_0403_));
 sky130_fd_sc_hd__a211o_1 _2750_ (.A1(_1311_),
    .A2(_1213_),
    .B1(_1449_),
    .C1(_0945_),
    .X(_0404_));
 sky130_fd_sc_hd__a211oi_1 _2751_ (.A1(_0786_),
    .A2(_0929_),
    .B1(_1174_),
    .C1(_1063_),
    .Y(_0405_));
 sky130_fd_sc_hd__a311oi_1 _2752_ (.A1(_0923_),
    .A2(_1392_),
    .A3(_1520_),
    .B1(_0405_),
    .C1(_1115_),
    .Y(_0406_));
 sky130_fd_sc_hd__a311o_1 _2753_ (.A1(_1278_),
    .A2(_0403_),
    .A3(_0404_),
    .B1(_0406_),
    .C1(_1193_),
    .X(_0407_));
 sky130_fd_sc_hd__a211o_1 _2754_ (.A1(_1219_),
    .A2(_1004_),
    .B1(_1084_),
    .C1(_1056_),
    .X(_0408_));
 sky130_fd_sc_hd__or2_1 _2755_ (.A(_0865_),
    .B(_1184_),
    .X(_0409_));
 sky130_fd_sc_hd__a221o_1 _2756_ (.A1(_0975_),
    .A2(_0976_),
    .B1(_1106_),
    .B2(_0802_),
    .C1(_0724_),
    .X(_0410_));
 sky130_fd_sc_hd__o311a_1 _2757_ (.A1(_1235_),
    .A2(_0966_),
    .A3(_1103_),
    .B1(_0410_),
    .C1(_0950_),
    .X(_0411_));
 sky130_fd_sc_hd__a311o_1 _2758_ (.A1(_1198_),
    .A2(_0408_),
    .A3(_0409_),
    .B1(_0411_),
    .C1(_0907_),
    .X(_0412_));
 sky130_fd_sc_hd__a21oi_1 _2759_ (.A1(_0407_),
    .A2(_0412_),
    .B1(_1039_),
    .Y(_0413_));
 sky130_fd_sc_hd__a311o_1 _2760_ (.A1(_0861_),
    .A2(_0402_),
    .A3(_1520_),
    .B1(_0413_),
    .C1(_0849_),
    .X(_0414_));
 sky130_fd_sc_hd__o311a_1 _2761_ (.A1(_1322_),
    .A2(_0388_),
    .A3(_0401_),
    .B1(_0414_),
    .C1(_0859_),
    .X(_0012_));
 sky130_fd_sc_hd__a21oi_2 _2762_ (.A1(_1219_),
    .A2(_1023_),
    .B1(_0762_),
    .Y(_0415_));
 sky130_fd_sc_hd__a211oi_4 _2763_ (.A1(_0734_),
    .A2(_0856_),
    .B1(_0415_),
    .C1(_0703_),
    .Y(_0416_));
 sky130_fd_sc_hd__nand2_1 _2764_ (.A(_0975_),
    .B(_1113_),
    .Y(_0417_));
 sky130_fd_sc_hd__o21a_1 _2765_ (.A1(_0805_),
    .A2(_0417_),
    .B1(_1095_),
    .X(_0418_));
 sky130_fd_sc_hd__o221a_1 _2766_ (.A1(_1299_),
    .A2(_0076_),
    .B1(_0418_),
    .B2(_0801_),
    .C1(_1115_),
    .X(_0419_));
 sky130_fd_sc_hd__a2111o_1 _2767_ (.A1(_0817_),
    .A2(_1077_),
    .B1(_1410_),
    .C1(_1050_),
    .D1(_0985_),
    .X(_0421_));
 sky130_fd_sc_hd__a21o_1 _2768_ (.A1(_0770_),
    .A2(_0340_),
    .B1(_1151_),
    .X(_0422_));
 sky130_fd_sc_hd__o21ai_1 _2769_ (.A1(_0764_),
    .A2(_0389_),
    .B1(_0964_),
    .Y(_0423_));
 sky130_fd_sc_hd__o311a_2 _2770_ (.A1(_0944_),
    .A2(_0940_),
    .A3(_1079_),
    .B1(_0423_),
    .C1(_0777_),
    .X(_0424_));
 sky130_fd_sc_hd__a311o_1 _2771_ (.A1(_1115_),
    .A2(_0421_),
    .A3(_0422_),
    .B1(_0424_),
    .C1(_0993_),
    .X(_0425_));
 sky130_fd_sc_hd__o311a_1 _2772_ (.A1(_0952_),
    .A2(_0416_),
    .A3(_0419_),
    .B1(_0425_),
    .C1(_0860_),
    .X(_0426_));
 sky130_fd_sc_hd__or3b_1 _2773_ (.A(_0964_),
    .B(_1064_),
    .C_N(_1475_),
    .X(_0427_));
 sky130_fd_sc_hd__o211a_1 _2774_ (.A1(_0900_),
    .A2(_0163_),
    .B1(_0427_),
    .C1(_0782_),
    .X(_0428_));
 sky130_fd_sc_hd__a21o_1 _2775_ (.A1(_0917_),
    .A2(_1152_),
    .B1(_1253_),
    .X(_0429_));
 sky130_fd_sc_hd__o311a_1 _2776_ (.A1(_1264_),
    .A2(_1190_),
    .A3(_1202_),
    .B1(_0429_),
    .C1(_1047_),
    .X(_0430_));
 sky130_fd_sc_hd__a211o_1 _2777_ (.A1(_0983_),
    .A2(_0948_),
    .B1(_1112_),
    .C1(_1140_),
    .X(_0431_));
 sky130_fd_sc_hd__a211o_1 _2778_ (.A1(_1124_),
    .A2(_1491_),
    .B1(_1524_),
    .C1(_0922_),
    .X(_0432_));
 sky130_fd_sc_hd__or3_1 _2779_ (.A(_0749_),
    .B(_0898_),
    .C(_1457_),
    .X(_0433_));
 sky130_fd_sc_hd__o211a_2 _2780_ (.A1(_1225_),
    .A2(_1330_),
    .B1(_0433_),
    .C1(_0777_),
    .X(_0434_));
 sky130_fd_sc_hd__a311o_1 _2781_ (.A1(_1047_),
    .A2(_0431_),
    .A3(_0432_),
    .B1(_0434_),
    .C1(_0993_),
    .X(_0435_));
 sky130_fd_sc_hd__o311a_1 _2782_ (.A1(_0952_),
    .A2(_0428_),
    .A3(_0430_),
    .B1(_0435_),
    .C1(_0645_),
    .X(_0436_));
 sky130_fd_sc_hd__o21ai_4 _2783_ (.A1(_0426_),
    .A2(_0436_),
    .B1(_0849_),
    .Y(_0437_));
 sky130_fd_sc_hd__o31ai_1 _2784_ (.A1(_1491_),
    .A2(_1016_),
    .A3(_1022_),
    .B1(_1211_),
    .Y(_0438_));
 sky130_fd_sc_hd__o311a_1 _2785_ (.A1(_1109_),
    .A2(_0940_),
    .A3(_0928_),
    .B1(_0438_),
    .C1(_1115_),
    .X(_0439_));
 sky130_fd_sc_hd__a211o_1 _2786_ (.A1(_0878_),
    .A2(_1173_),
    .B1(_1466_),
    .C1(_0922_),
    .X(_0440_));
 sky130_fd_sc_hd__o211a_1 _2787_ (.A1(_0075_),
    .A2(_0158_),
    .B1(_0440_),
    .C1(_0782_),
    .X(_0442_));
 sky130_fd_sc_hd__or3b_1 _2788_ (.A(_0345_),
    .B(_0724_),
    .C_N(_1098_),
    .X(_0443_));
 sky130_fd_sc_hd__nor2_1 _2789_ (.A(_1391_),
    .B(_1078_),
    .Y(_0444_));
 sky130_fd_sc_hd__or3_1 _2790_ (.A(_0910_),
    .B(_1043_),
    .C(_0444_),
    .X(_0445_));
 sky130_fd_sc_hd__a311o_1 _2791_ (.A1(_0825_),
    .A2(_1015_),
    .A3(_0946_),
    .B1(_1236_),
    .C1(_0749_),
    .X(_0446_));
 sky130_fd_sc_hd__o311a_1 _2792_ (.A1(_0944_),
    .A2(_0821_),
    .A3(_0146_),
    .B1(_0446_),
    .C1(_0838_),
    .X(_0447_));
 sky130_fd_sc_hd__a311o_1 _2793_ (.A1(_0978_),
    .A2(_0443_),
    .A3(_0445_),
    .B1(_0447_),
    .C1(_0842_),
    .X(_0448_));
 sky130_fd_sc_hd__o311a_2 _2794_ (.A1(_0667_),
    .A2(_0439_),
    .A3(_0442_),
    .B1(_0448_),
    .C1(_1036_),
    .X(_0449_));
 sky130_fd_sc_hd__a21oi_4 _2795_ (.A1(_0881_),
    .A2(_0797_),
    .B1(_0769_),
    .Y(_0450_));
 sky130_fd_sc_hd__o31a_1 _2796_ (.A1(_0787_),
    .A2(_0901_),
    .A3(_0450_),
    .B1(_0860_),
    .X(_0451_));
 sky130_fd_sc_hd__o21ai_1 _2797_ (.A1(_0449_),
    .A2(_0451_),
    .B1(_0863_),
    .Y(_0453_));
 sky130_fd_sc_hd__and3_1 _2798_ (.A(net66),
    .B(_0437_),
    .C(net71),
    .X(_0454_));
 sky130_fd_sc_hd__buf_1 _2799_ (.A(net72),
    .X(_0013_));
 sky130_fd_sc_hd__o211ai_1 _2800_ (.A1(_1343_),
    .A2(_1020_),
    .B1(_1055_),
    .C1(_0811_),
    .Y(_0455_));
 sky130_fd_sc_hd__o311a_1 _2801_ (.A1(_1274_),
    .A2(_1045_),
    .A3(_1094_),
    .B1(_0455_),
    .C1(_0935_),
    .X(_0456_));
 sky130_fd_sc_hd__a311o_1 _2802_ (.A1(_1199_),
    .A2(_1219_),
    .A3(_0947_),
    .B1(_1172_),
    .C1(_0957_),
    .X(_0457_));
 sky130_fd_sc_hd__o311a_1 _2803_ (.A1(_1345_),
    .A2(_0855_),
    .A3(_1213_),
    .B1(_0457_),
    .C1(_1287_),
    .X(_0458_));
 sky130_fd_sc_hd__or3_1 _2804_ (.A(_1164_),
    .B(_0456_),
    .C(_0458_),
    .X(_0459_));
 sky130_fd_sc_hd__nand2_1 _2805_ (.A(_1274_),
    .B(_0919_),
    .Y(_0460_));
 sky130_fd_sc_hd__or3_1 _2806_ (.A(_0873_),
    .B(_1491_),
    .C(_1463_),
    .X(_0461_));
 sky130_fd_sc_hd__o211a_1 _2807_ (.A1(_0460_),
    .A2(_0344_),
    .B1(_0461_),
    .C1(_1285_),
    .X(_0463_));
 sky130_fd_sc_hd__or3_1 _2808_ (.A(_1491_),
    .B(_1016_),
    .C(_0353_),
    .X(_0464_));
 sky130_fd_sc_hd__o311a_1 _2809_ (.A1(_1403_),
    .A2(_1119_),
    .A3(_0273_),
    .B1(_0464_),
    .C1(_1308_),
    .X(_0465_));
 sky130_fd_sc_hd__o31a_1 _2810_ (.A1(_1298_),
    .A2(_0463_),
    .A3(_0465_),
    .B1(_1039_),
    .X(_0466_));
 sky130_fd_sc_hd__and3_2 _2811_ (.A(_0769_),
    .B(_0999_),
    .C(_0851_),
    .X(_0467_));
 sky130_fd_sc_hd__or3_1 _2812_ (.A(_0936_),
    .B(_0888_),
    .C(_0124_),
    .X(_0468_));
 sky130_fd_sc_hd__o311a_1 _2813_ (.A1(_1348_),
    .A2(_1516_),
    .A3(_0467_),
    .B1(_0468_),
    .C1(_1285_),
    .X(_0469_));
 sky130_fd_sc_hd__a211o_1 _2814_ (.A1(_1347_),
    .A2(_0973_),
    .B1(_0214_),
    .C1(_0923_),
    .X(_0470_));
 sky130_fd_sc_hd__o311a_1 _2815_ (.A1(_1281_),
    .A2(_0990_),
    .A3(_1470_),
    .B1(_0470_),
    .C1(_1308_),
    .X(_0471_));
 sky130_fd_sc_hd__a21o_1 _2816_ (.A1(_0916_),
    .A2(_1077_),
    .B1(_1023_),
    .X(_0472_));
 sky130_fd_sc_hd__nand2_1 _2817_ (.A(_0936_),
    .B(_1399_),
    .Y(_0474_));
 sky130_fd_sc_hd__xnor2_1 _2818_ (.A(_0472_),
    .B(_0474_),
    .Y(_0475_));
 sky130_fd_sc_hd__a211o_1 _2819_ (.A1(_0878_),
    .A2(_1213_),
    .B1(_0450_),
    .C1(_1140_),
    .X(_0476_));
 sky130_fd_sc_hd__o311a_1 _2820_ (.A1(_0751_),
    .A2(_1418_),
    .A3(_1449_),
    .B1(_0476_),
    .C1(_0782_),
    .X(_0477_));
 sky130_fd_sc_hd__a211o_1 _2821_ (.A1(_1342_),
    .A2(_0475_),
    .B1(_0477_),
    .C1(_0952_),
    .X(_0478_));
 sky130_fd_sc_hd__o311a_1 _2822_ (.A1(_0673_),
    .A2(_0469_),
    .A3(_0471_),
    .B1(_0478_),
    .C1(_1396_),
    .X(_0479_));
 sky130_fd_sc_hd__a21oi_1 _2823_ (.A1(_0459_),
    .A2(_0466_),
    .B1(_0479_),
    .Y(_0480_));
 sky130_fd_sc_hd__a221o_1 _2824_ (.A1(_1000_),
    .A2(_1229_),
    .B1(_0819_),
    .B2(_1199_),
    .C1(_1109_),
    .X(_0481_));
 sky130_fd_sc_hd__o311a_1 _2825_ (.A1(_1348_),
    .A2(_1044_),
    .A3(_1487_),
    .B1(_0481_),
    .C1(_0935_),
    .X(_0482_));
 sky130_fd_sc_hd__or3_1 _2826_ (.A(_0873_),
    .B(_1292_),
    .C(_0266_),
    .X(_0483_));
 sky130_fd_sc_hd__o311a_1 _2827_ (.A1(_1345_),
    .A2(_0813_),
    .A3(_1466_),
    .B1(_0483_),
    .C1(_1287_),
    .X(_0485_));
 sky130_fd_sc_hd__nor2_1 _2828_ (.A(_1347_),
    .B(_1073_),
    .Y(_0486_));
 sky130_fd_sc_hd__a211o_1 _2829_ (.A1(_1053_),
    .A2(_1073_),
    .B1(_1165_),
    .C1(_0827_),
    .X(_0487_));
 sky130_fd_sc_hd__o311a_1 _2830_ (.A1(_0752_),
    .A2(_1182_),
    .A3(_0486_),
    .B1(_0487_),
    .C1(_1342_),
    .X(_0488_));
 sky130_fd_sc_hd__a311o_1 _2831_ (.A1(_1343_),
    .A2(_1019_),
    .A3(_0971_),
    .B1(_1189_),
    .C1(_0911_),
    .X(_0489_));
 sky130_fd_sc_hd__a311o_1 _2832_ (.A1(_1232_),
    .A2(_1367_),
    .A3(_0867_),
    .B1(_1152_),
    .C1(_0801_),
    .X(_0490_));
 sky130_fd_sc_hd__a31o_1 _2833_ (.A1(_1356_),
    .A2(_0489_),
    .A3(_0490_),
    .B1(_0952_),
    .X(_0491_));
 sky130_fd_sc_hd__o32a_1 _2834_ (.A1(_1164_),
    .A2(_0482_),
    .A3(_0485_),
    .B1(_0488_),
    .B2(_0491_),
    .X(_0492_));
 sky130_fd_sc_hd__a211o_1 _2835_ (.A1(_0917_),
    .A2(_1379_),
    .B1(_0270_),
    .C1(_1161_),
    .X(_0493_));
 sky130_fd_sc_hd__o211ai_1 _2836_ (.A1(_1365_),
    .A2(_0492_),
    .B1(_0493_),
    .C1(_1322_),
    .Y(_0494_));
 sky130_fd_sc_hd__o211a_1 _2837_ (.A1(_1322_),
    .A2(_0480_),
    .B1(_0494_),
    .C1(_1242_),
    .X(_0014_));
 sky130_fd_sc_hd__a211o_1 _2838_ (.A1(_1206_),
    .A2(_0172_),
    .B1(_1457_),
    .C1(_1281_),
    .X(_0496_));
 sky130_fd_sc_hd__a21o_1 _2839_ (.A1(_1055_),
    .A2(_1359_),
    .B1(_0752_),
    .X(_0497_));
 sky130_fd_sc_hd__or3_1 _2840_ (.A(_1063_),
    .B(_1249_),
    .C(_0467_),
    .X(_0498_));
 sky130_fd_sc_hd__o211a_1 _2841_ (.A1(_1252_),
    .A2(_0316_),
    .B1(_0498_),
    .C1(_0935_),
    .X(_0499_));
 sky130_fd_sc_hd__a311oi_1 _2842_ (.A1(_0706_),
    .A2(_0496_),
    .A3(_0497_),
    .B1(_0499_),
    .C1(_1243_),
    .Y(_0500_));
 sky130_fd_sc_hd__o22a_1 _2843_ (.A1(_0801_),
    .A2(_0977_),
    .B1(_1137_),
    .B2(_1043_),
    .X(_0501_));
 sky130_fd_sc_hd__a31o_1 _2844_ (.A1(_0828_),
    .A2(_1244_),
    .A3(_1084_),
    .B1(_0501_),
    .X(_0502_));
 sky130_fd_sc_hd__a211o_1 _2845_ (.A1(_0721_),
    .A2(_0739_),
    .B1(_1106_),
    .C1(_1165_),
    .X(_0503_));
 sky130_fd_sc_hd__a211o_1 _2846_ (.A1(_1232_),
    .A2(_1127_),
    .B1(_1410_),
    .C1(_1261_),
    .X(_0504_));
 sky130_fd_sc_hd__a31o_1 _2847_ (.A1(_0783_),
    .A2(_0503_),
    .A3(_0504_),
    .B1(_1318_),
    .X(_0506_));
 sky130_fd_sc_hd__a21oi_1 _2848_ (.A1(_0706_),
    .A2(_0502_),
    .B1(_0506_),
    .Y(_0507_));
 sky130_fd_sc_hd__or3b_1 _2849_ (.A(_0911_),
    .B(_0827_),
    .C_N(_1359_),
    .X(_0508_));
 sky130_fd_sc_hd__a21o_1 _2850_ (.A1(_0917_),
    .A2(_0807_),
    .B1(_1389_),
    .X(_0509_));
 sky130_fd_sc_hd__nand3_1 _2851_ (.A(_1250_),
    .B(_0508_),
    .C(_0509_),
    .Y(_0510_));
 sky130_fd_sc_hd__o21a_1 _2852_ (.A1(_0827_),
    .A2(_0105_),
    .B1(_1180_),
    .X(_0511_));
 sky130_fd_sc_hd__a311o_1 _2853_ (.A1(_0734_),
    .A2(_1146_),
    .A3(_1167_),
    .B1(_0511_),
    .C1(_1178_),
    .X(_0512_));
 sky130_fd_sc_hd__o21a_1 _2854_ (.A1(_1059_),
    .A2(_0444_),
    .B1(_0944_),
    .X(_0513_));
 sky130_fd_sc_hd__a311o_1 _2855_ (.A1(_1056_),
    .A2(_0871_),
    .A3(_1055_),
    .B1(_0513_),
    .C1(_0694_),
    .X(_0514_));
 sky130_fd_sc_hd__nor3_1 _2856_ (.A(_1060_),
    .B(_0815_),
    .C(_1118_),
    .Y(_0515_));
 sky130_fd_sc_hd__a311o_1 _2857_ (.A1(_0936_),
    .A2(_0390_),
    .A3(_0186_),
    .B1(_0515_),
    .C1(_0934_),
    .X(_0517_));
 sky130_fd_sc_hd__a31o_1 _2858_ (.A1(_0907_),
    .A2(_0514_),
    .A3(_0517_),
    .B1(_0860_),
    .X(_0518_));
 sky130_fd_sc_hd__a31o_1 _2859_ (.A1(_1298_),
    .A2(_0510_),
    .A3(_0512_),
    .B1(_0518_),
    .X(_0519_));
 sky130_fd_sc_hd__o31a_1 _2860_ (.A1(_1396_),
    .A2(_0500_),
    .A3(_0507_),
    .B1(_0519_),
    .X(_0520_));
 sky130_fd_sc_hd__or3b_1 _2861_ (.A(_1400_),
    .B(_0725_),
    .C_N(_0722_),
    .X(_0521_));
 sky130_fd_sc_hd__o311a_1 _2862_ (.A1(_1345_),
    .A2(_0270_),
    .A3(_0303_),
    .B1(_0521_),
    .C1(_0779_),
    .X(_0522_));
 sky130_fd_sc_hd__or3b_1 _2863_ (.A(_1467_),
    .B(_0875_),
    .C_N(_1160_),
    .X(_0523_));
 sky130_fd_sc_hd__a211o_1 _2864_ (.A1(_0803_),
    .A2(_1099_),
    .B1(_1142_),
    .C1(_1040_),
    .X(_0524_));
 sky130_fd_sc_hd__and3_2 _2865_ (.A(_1278_),
    .B(_0523_),
    .C(_0524_),
    .X(_0525_));
 sky130_fd_sc_hd__o21ai_1 _2866_ (.A1(_0522_),
    .A2(_0525_),
    .B1(_0673_),
    .Y(_0526_));
 sky130_fd_sc_hd__mux2_1 _2867_ (.A0(_0940_),
    .A1(_1487_),
    .S(_0873_),
    .X(_0528_));
 sky130_fd_sc_hd__o21a_1 _2868_ (.A1(_0221_),
    .A2(_0528_),
    .B1(_1356_),
    .X(_0529_));
 sky130_fd_sc_hd__o221ai_2 _2869_ (.A1(_1343_),
    .A2(_0996_),
    .B1(_0940_),
    .B2(_1261_),
    .C1(_1329_),
    .Y(_0530_));
 sky130_fd_sc_hd__o311a_1 _2870_ (.A1(_1403_),
    .A2(_1379_),
    .A3(_0124_),
    .B1(_0530_),
    .C1(_1308_),
    .X(_0531_));
 sky130_fd_sc_hd__o21ai_1 _2871_ (.A1(_0529_),
    .A2(_0531_),
    .B1(_1243_),
    .Y(_0532_));
 sky130_fd_sc_hd__o211a_1 _2872_ (.A1(_1124_),
    .A2(_0880_),
    .B1(_1532_),
    .C1(_1039_),
    .X(_0533_));
 sky130_fd_sc_hd__a311o_1 _2873_ (.A1(_0655_),
    .A2(_0526_),
    .A3(_0532_),
    .B1(_0533_),
    .C1(_0849_),
    .X(_0534_));
 sky130_fd_sc_hd__o211a_1 _2874_ (.A1(_1322_),
    .A2(_0520_),
    .B1(_0534_),
    .C1(_1242_),
    .X(_0016_));
 sky130_fd_sc_hd__or3_1 _2875_ (.A(_0724_),
    .B(_0747_),
    .C(_1277_),
    .X(_0535_));
 sky130_fd_sc_hd__o311a_1 _2876_ (.A1(_1109_),
    .A2(_1432_),
    .A3(_0467_),
    .B1(_0535_),
    .C1(_0978_),
    .X(_0536_));
 sky130_fd_sc_hd__a211o_1 _2877_ (.A1(_1229_),
    .A2(_1399_),
    .B1(_1380_),
    .C1(_1083_),
    .X(_0538_));
 sky130_fd_sc_hd__o311a_2 _2878_ (.A1(_1040_),
    .A2(_1059_),
    .A3(_0289_),
    .B1(_0538_),
    .C1(_1047_),
    .X(_0539_));
 sky130_fd_sc_hd__a221o_1 _2879_ (.A1(_1078_),
    .A2(_1221_),
    .B1(_0959_),
    .B2(_0931_),
    .C1(_0749_),
    .X(_0540_));
 sky130_fd_sc_hd__o311a_1 _2880_ (.A1(_0964_),
    .A2(_1026_),
    .A3(_1168_),
    .B1(_0540_),
    .C1(_0838_),
    .X(_0541_));
 sky130_fd_sc_hd__o21ai_1 _2881_ (.A1(_0767_),
    .A2(_0931_),
    .B1(_1028_),
    .Y(_0542_));
 sky130_fd_sc_hd__a21oi_1 _2882_ (.A1(_1187_),
    .A2(_0542_),
    .B1(_0694_),
    .Y(_0543_));
 sky130_fd_sc_hd__or3_1 _2883_ (.A(_0661_),
    .B(_0541_),
    .C(_0543_),
    .X(_0544_));
 sky130_fd_sc_hd__o311a_1 _2884_ (.A1(_1193_),
    .A2(_0536_),
    .A3(_0539_),
    .B1(_0544_),
    .C1(_0860_),
    .X(_0545_));
 sky130_fd_sc_hd__a2bb2o_1 _2885_ (.A1_N(_0970_),
    .A2_N(_1213_),
    .B1(_0744_),
    .B2(_0739_),
    .X(_0546_));
 sky130_fd_sc_hd__a211o_1 _2886_ (.A1(_0786_),
    .A2(_0868_),
    .B1(_1202_),
    .C1(_1140_),
    .X(_0547_));
 sky130_fd_sc_hd__o211a_1 _2887_ (.A1(_0923_),
    .A2(_0546_),
    .B1(_0547_),
    .C1(_1047_),
    .X(_0549_));
 sky130_fd_sc_hd__a221o_1 _2888_ (.A1(_1019_),
    .A2(_1043_),
    .B1(_1206_),
    .B2(_0172_),
    .C1(_1140_),
    .X(_0550_));
 sky130_fd_sc_hd__o311a_1 _2889_ (.A1(_0801_),
    .A2(_0890_),
    .A3(_1150_),
    .B1(_0550_),
    .C1(_0782_),
    .X(_0551_));
 sky130_fd_sc_hd__o21ai_1 _2890_ (.A1(_0724_),
    .A2(_0899_),
    .B1(_1219_),
    .Y(_0552_));
 sky130_fd_sc_hd__a32o_1 _2891_ (.A1(_1089_),
    .A2(_1083_),
    .A3(_0770_),
    .B1(_0552_),
    .B2(_1124_),
    .X(_0553_));
 sky130_fd_sc_hd__a21oi_1 _2892_ (.A1(_0772_),
    .A2(_0712_),
    .B1(_0826_),
    .Y(_0554_));
 sky130_fd_sc_hd__or4_1 _2893_ (.A(_0723_),
    .B(_0890_),
    .C(_1168_),
    .D(_0554_),
    .X(_0555_));
 sky130_fd_sc_hd__o311a_1 _2894_ (.A1(_1060_),
    .A2(_1422_),
    .A3(_0154_),
    .B1(_0555_),
    .C1(_0914_),
    .X(_0556_));
 sky130_fd_sc_hd__a211o_1 _2895_ (.A1(_0839_),
    .A2(_0553_),
    .B1(_0556_),
    .C1(_0842_),
    .X(_0557_));
 sky130_fd_sc_hd__o311a_1 _2896_ (.A1(_1318_),
    .A2(_0549_),
    .A3(_0551_),
    .B1(_0557_),
    .C1(_1036_),
    .X(_0558_));
 sky130_fd_sc_hd__o21ai_4 _2897_ (.A1(_0545_),
    .A2(_0558_),
    .B1(_0849_),
    .Y(_0560_));
 sky130_fd_sc_hd__a21o_1 _2898_ (.A1(_0785_),
    .A2(_0380_),
    .B1(_0749_),
    .X(_0561_));
 sky130_fd_sc_hd__o32a_1 _2899_ (.A1(_0964_),
    .A2(_0941_),
    .A3(_1230_),
    .B1(_0561_),
    .B2(_0913_),
    .X(_0562_));
 sky130_fd_sc_hd__o31a_1 _2900_ (.A1(_0944_),
    .A2(_0948_),
    .A3(_1433_),
    .B1(_0777_),
    .X(_0563_));
 sky130_fd_sc_hd__or2b_1 _2901_ (.A(_0561_),
    .B_N(_1329_),
    .X(_0564_));
 sky130_fd_sc_hd__a2bb2o_1 _2902_ (.A1_N(_0934_),
    .A2_N(_0562_),
    .B1(_0563_),
    .B2(_0564_),
    .X(_0565_));
 sky130_fd_sc_hd__a221o_1 _2903_ (.A1(_0721_),
    .A2(_0739_),
    .B1(_1072_),
    .B2(_1159_),
    .C1(_0956_),
    .X(_0566_));
 sky130_fd_sc_hd__a21o_1 _2904_ (.A1(_0824_),
    .A2(_1106_),
    .B1(_0358_),
    .X(_0567_));
 sky130_fd_sc_hd__a221o_1 _2905_ (.A1(_0802_),
    .A2(_1105_),
    .B1(_1324_),
    .B2(_0892_),
    .C1(_0834_),
    .X(_0568_));
 sky130_fd_sc_hd__o311a_1 _2906_ (.A1(_0956_),
    .A2(_0744_),
    .A3(_1172_),
    .B1(_0568_),
    .C1(_0838_),
    .X(_0569_));
 sky130_fd_sc_hd__a311o_1 _2907_ (.A1(_0778_),
    .A2(_0566_),
    .A3(_0567_),
    .B1(_0569_),
    .C1(_0841_),
    .X(_0571_));
 sky130_fd_sc_hd__o21ai_2 _2908_ (.A1(_1318_),
    .A2(_0565_),
    .B1(_0571_),
    .Y(_0572_));
 sky130_fd_sc_hd__nor2_1 _2909_ (.A(_1036_),
    .B(_0075_),
    .Y(_0573_));
 sky130_fd_sc_hd__a221o_1 _2910_ (.A1(_0645_),
    .A2(_0572_),
    .B1(_0573_),
    .B2(_1497_),
    .C1(_0848_),
    .X(_0574_));
 sky130_fd_sc_hd__and3_1 _2911_ (.A(net66),
    .B(_0560_),
    .C(_0574_),
    .X(_0575_));
 sky130_fd_sc_hd__buf_1 _2912_ (.A(_0575_),
    .X(_0017_));
 sky130_fd_sc_hd__nor2_1 _2913_ (.A(_1125_),
    .B(_0124_),
    .Y(_0576_));
 sky130_fd_sc_hd__o21ai_1 _2914_ (.A1(_1111_),
    .A2(_0209_),
    .B1(_1049_),
    .Y(_0577_));
 sky130_fd_sc_hd__o311ai_4 _2915_ (.A1(_1235_),
    .A2(_1141_),
    .A3(_1500_),
    .B1(_0577_),
    .C1(_0694_),
    .Y(_0578_));
 sky130_fd_sc_hd__o21ai_1 _2916_ (.A1(_0855_),
    .A2(_0331_),
    .B1(_0985_),
    .Y(_0579_));
 sky130_fd_sc_hd__o21ai_1 _2917_ (.A1(_0928_),
    .A2(_0450_),
    .B1(_0800_),
    .Y(_0581_));
 sky130_fd_sc_hd__a21o_1 _2918_ (.A1(_0579_),
    .A2(_0581_),
    .B1(_0694_),
    .X(_0582_));
 sky130_fd_sc_hd__o21ai_2 _2919_ (.A1(_1099_),
    .A2(_1407_),
    .B1(_0749_),
    .Y(_0583_));
 sky130_fd_sc_hd__o311a_1 _2920_ (.A1(_0799_),
    .A2(_1466_),
    .A3(_0075_),
    .B1(_0583_),
    .C1(_0776_),
    .X(_0584_));
 sky130_fd_sc_hd__or3_1 _2921_ (.A(_0833_),
    .B(_0768_),
    .C(_0965_),
    .X(_0585_));
 sky130_fd_sc_hd__o21ai_1 _2922_ (.A1(_1265_),
    .A2(_1334_),
    .B1(_0984_),
    .Y(_0586_));
 sky130_fd_sc_hd__and3_1 _2923_ (.A(_0685_),
    .B(_0585_),
    .C(_0586_),
    .X(_0587_));
 sky130_fd_sc_hd__o21a_1 _2924_ (.A1(_0584_),
    .A2(_0587_),
    .B1(_0841_),
    .X(_0588_));
 sky130_fd_sc_hd__a31o_1 _2925_ (.A1(_0907_),
    .A2(_0578_),
    .A3(_0582_),
    .B1(_0588_),
    .X(_0589_));
 sky130_fd_sc_hd__and3_2 _2926_ (.A(_0926_),
    .B(_0713_),
    .C(_0999_),
    .X(_0590_));
 sky130_fd_sc_hd__a211o_1 _2927_ (.A1(_0825_),
    .A2(_1077_),
    .B1(_0137_),
    .C1(_0749_),
    .X(_0592_));
 sky130_fd_sc_hd__o311a_1 _2928_ (.A1(_0964_),
    .A2(_1276_),
    .A3(_0590_),
    .B1(_0592_),
    .C1(_0777_),
    .X(_0593_));
 sky130_fd_sc_hd__and3_1 _2929_ (.A(_0716_),
    .B(_0924_),
    .C(_0959_),
    .X(_0594_));
 sky130_fd_sc_hd__o21ai_4 _2930_ (.A1(_1432_),
    .A2(_0594_),
    .B1(_1028_),
    .Y(_0595_));
 sky130_fd_sc_hd__a211o_1 _2931_ (.A1(_1117_),
    .A2(_0896_),
    .B1(_0887_),
    .C1(_0864_),
    .X(_0596_));
 sky130_fd_sc_hd__a21oi_1 _2932_ (.A1(_0595_),
    .A2(_0596_),
    .B1(_0914_),
    .Y(_0597_));
 sky130_fd_sc_hd__nor2_1 _2933_ (.A(_0593_),
    .B(_0597_),
    .Y(_0598_));
 sky130_fd_sc_hd__o211ai_1 _2934_ (.A1(_1127_),
    .A2(_1422_),
    .B1(_0910_),
    .C1(_1232_),
    .Y(_0599_));
 sky130_fd_sc_hd__o21ai_1 _2935_ (.A1(_0771_),
    .A2(_0389_),
    .B1(_0956_),
    .Y(_0600_));
 sky130_fd_sc_hd__o211a_1 _2936_ (.A1(_0745_),
    .A2(_1073_),
    .B1(_0257_),
    .C1(_0723_),
    .X(_0601_));
 sky130_fd_sc_hd__o221a_1 _2937_ (.A1(_0791_),
    .A2(_0805_),
    .B1(_1392_),
    .B2(_1078_),
    .C1(_0833_),
    .X(_0603_));
 sky130_fd_sc_hd__o21a_1 _2938_ (.A1(_0601_),
    .A2(_0603_),
    .B1(_0776_),
    .X(_0604_));
 sky130_fd_sc_hd__a311o_2 _2939_ (.A1(_0838_),
    .A2(_0599_),
    .A3(_0600_),
    .B1(_0604_),
    .C1(_0841_),
    .X(_0605_));
 sky130_fd_sc_hd__o21a_1 _2940_ (.A1(_0907_),
    .A2(_0598_),
    .B1(_0605_),
    .X(_0606_));
 sky130_fd_sc_hd__a21o_1 _2941_ (.A1(_0264_),
    .A2(_0093_),
    .B1(_0755_),
    .X(_0607_));
 sky130_fd_sc_hd__or3_4 _2942_ (.A(_0910_),
    .B(_0948_),
    .C(_0913_),
    .X(_0608_));
 sky130_fd_sc_hd__a21oi_1 _2943_ (.A1(_0607_),
    .A2(_0608_),
    .B1(_0782_),
    .Y(_0609_));
 sky130_fd_sc_hd__a211o_1 _2944_ (.A1(_1013_),
    .A2(_1106_),
    .B1(_0303_),
    .C1(_0944_),
    .X(_0610_));
 sky130_fd_sc_hd__o311a_1 _2945_ (.A1(_0875_),
    .A2(_1206_),
    .A3(_1130_),
    .B1(_0610_),
    .C1(_0934_),
    .X(_0611_));
 sky130_fd_sc_hd__a221o_1 _2946_ (.A1(_1136_),
    .A2(_1031_),
    .B1(_0983_),
    .B2(_0931_),
    .C1(_0956_),
    .X(_0612_));
 sky130_fd_sc_hd__a211o_1 _2947_ (.A1(_1011_),
    .A2(_0787_),
    .B1(_1354_),
    .C1(_1028_),
    .X(_0614_));
 sky130_fd_sc_hd__or3_1 _2948_ (.A(_0834_),
    .B(_1247_),
    .C(_1306_),
    .X(_0615_));
 sky130_fd_sc_hd__or3_1 _2949_ (.A(_0723_),
    .B(_0764_),
    .C(_0888_),
    .X(_0616_));
 sky130_fd_sc_hd__a31o_2 _2950_ (.A1(_0685_),
    .A2(_0615_),
    .A3(_0616_),
    .B1(_0661_),
    .X(_0617_));
 sky130_fd_sc_hd__a31o_1 _2951_ (.A1(_0778_),
    .A2(_0612_),
    .A3(_0614_),
    .B1(_0617_),
    .X(_0618_));
 sky130_fd_sc_hd__o31ai_1 _2952_ (.A1(_1193_),
    .A2(_0609_),
    .A3(_0611_),
    .B1(_0618_),
    .Y(_0619_));
 sky130_fd_sc_hd__mux4_1 _2953_ (.A0(_0576_),
    .A1(_0589_),
    .A2(_0606_),
    .A3(_0619_),
    .S0(_1036_),
    .S1(_0848_),
    .X(_0620_));
 sky130_fd_sc_hd__and2_1 _2954_ (.A(_0859_),
    .B(_0620_),
    .X(_0621_));
 sky130_fd_sc_hd__clkbuf_1 _2955_ (.A(_0621_),
    .X(_0018_));
 sky130_fd_sc_hd__o21ai_1 _2956_ (.A1(_0744_),
    .A2(_1130_),
    .B1(_1261_),
    .Y(_0622_));
 sky130_fd_sc_hd__a21o_1 _2957_ (.A1(_0579_),
    .A2(_0622_),
    .B1(_0703_),
    .X(_0624_));
 sky130_fd_sc_hd__a21o_1 _2958_ (.A1(_0578_),
    .A2(_0624_),
    .B1(_0843_),
    .X(_0625_));
 sky130_fd_sc_hd__o21ai_1 _2959_ (.A1(_1182_),
    .A2(_1224_),
    .B1(_1244_),
    .Y(_0626_));
 sky130_fd_sc_hd__a21oi_1 _2960_ (.A1(_0771_),
    .A2(_1146_),
    .B1(_0744_),
    .Y(_0627_));
 sky130_fd_sc_hd__o211a_1 _2961_ (.A1(_0811_),
    .A2(_0627_),
    .B1(_0585_),
    .C1(_0839_),
    .X(_0628_));
 sky130_fd_sc_hd__a311o_1 _2962_ (.A1(_1250_),
    .A2(_0583_),
    .A3(_0626_),
    .B1(_0628_),
    .C1(_1164_),
    .X(_0629_));
 sky130_fd_sc_hd__o211a_1 _2963_ (.A1(_1396_),
    .A2(_1181_),
    .B1(_0625_),
    .C1(_0629_),
    .X(_0630_));
 sky130_fd_sc_hd__a21oi_1 _2964_ (.A1(_0625_),
    .A2(_0629_),
    .B1(_0655_),
    .Y(_0631_));
 sky130_fd_sc_hd__a211o_1 _2965_ (.A1(_1367_),
    .A2(_1254_),
    .B1(_0137_),
    .C1(_0957_),
    .X(_0632_));
 sky130_fd_sc_hd__o311a_1 _2966_ (.A1(_1335_),
    .A2(_0721_),
    .A3(_0590_),
    .B1(_0632_),
    .C1(_0935_),
    .X(_0633_));
 sky130_fd_sc_hd__a21o_1 _2967_ (.A1(_0110_),
    .A2(_0186_),
    .B1(_1256_),
    .X(_0635_));
 sky130_fd_sc_hd__a21oi_1 _2968_ (.A1(_0595_),
    .A2(_0635_),
    .B1(_0783_),
    .Y(_0636_));
 sky130_fd_sc_hd__o21ai_1 _2969_ (.A1(_0633_),
    .A2(_0636_),
    .B1(_1243_),
    .Y(_0637_));
 sky130_fd_sc_hd__a21oi_1 _2970_ (.A1(_0605_),
    .A2(_0637_),
    .B1(_1396_),
    .Y(_0638_));
 sky130_fd_sc_hd__a21oi_1 _2971_ (.A1(_0824_),
    .A2(_0807_),
    .B1(_0130_),
    .Y(_0639_));
 sky130_fd_sc_hd__o21ai_1 _2972_ (.A1(_1291_),
    .A2(_0639_),
    .B1(_0608_),
    .Y(_0640_));
 sky130_fd_sc_hd__nand2_1 _2973_ (.A(_1211_),
    .B(_1120_),
    .Y(_0641_));
 sky130_fd_sc_hd__a211o_1 _2974_ (.A1(_1013_),
    .A2(_1314_),
    .B1(_0303_),
    .C1(_0985_),
    .X(_0642_));
 sky130_fd_sc_hd__o211a_1 _2975_ (.A1(_0807_),
    .A2(_0641_),
    .B1(_0642_),
    .C1(_0778_),
    .X(_0643_));
 sky130_fd_sc_hd__a211o_1 _2976_ (.A1(_1310_),
    .A2(_0640_),
    .B1(_0643_),
    .C1(_0952_),
    .X(_0644_));
 sky130_fd_sc_hd__a211o_1 _2977_ (.A1(_1347_),
    .A2(_0787_),
    .B1(_1206_),
    .C1(_0911_),
    .X(_0646_));
 sky130_fd_sc_hd__a211o_1 _2978_ (.A1(_0983_),
    .A2(_0931_),
    .B1(_1300_),
    .C1(_0923_),
    .X(_0647_));
 sky130_fd_sc_hd__a31o_1 _2979_ (.A1(_1356_),
    .A2(_0646_),
    .A3(_0647_),
    .B1(_0617_),
    .X(_0648_));
 sky130_fd_sc_hd__and3_1 _2980_ (.A(_1161_),
    .B(_0644_),
    .C(_0648_),
    .X(_0649_));
 sky130_fd_sc_hd__o21ai_1 _2981_ (.A1(_0638_),
    .A2(_0649_),
    .B1(_1197_),
    .Y(_0650_));
 sky130_fd_sc_hd__o311a_1 _2982_ (.A1(_1197_),
    .A2(_0630_),
    .A3(_0631_),
    .B1(_0859_),
    .C1(_0650_),
    .X(_0020_));
 sky130_fd_sc_hd__or4_1 _2983_ (.A(net8),
    .B(net9),
    .C(net10),
    .D(net85),
    .X(_0651_));
 sky130_fd_sc_hd__or4b_1 _2984_ (.A(net6),
    .B(net4),
    .C(net7),
    .D_N(net5),
    .X(_0652_));
 sky130_fd_sc_hd__nor4_1 _2985_ (.A(net18),
    .B(_0420_),
    .C(_0651_),
    .D(_0652_),
    .Y(_0653_));
 sky130_fd_sc_hd__buf_2 _2986_ (.A(_0653_),
    .X(_0654_));
 sky130_fd_sc_hd__or4_1 _2987_ (.A(net6),
    .B(net4),
    .C(net7),
    .D(net5),
    .X(_0656_));
 sky130_fd_sc_hd__or2_1 _2988_ (.A(_0651_),
    .B(_0656_),
    .X(_0657_));
 sky130_fd_sc_hd__nor3_1 _2989_ (.A(net18),
    .B(_0420_),
    .C(_0657_),
    .Y(_0658_));
 sky130_fd_sc_hd__a22o_1 _2990_ (.A1(\weights_inst.data_out[0] ),
    .A2(_0654_),
    .B1(net53),
    .B2(\fsm_inst.cnn_en ),
    .X(net20));
 sky130_fd_sc_hd__a22o_1 _2991_ (.A1(\weights_inst.data_out[1] ),
    .A2(_0654_),
    .B1(net53),
    .B2(\fsm_inst.batch_norm_en ),
    .X(net31));
 sky130_fd_sc_hd__a22o_1 _2992_ (.A1(\weights_inst.data_out[2] ),
    .A2(_0654_),
    .B1(_0658_),
    .B2(\fsm_inst.done ),
    .X(net42));
 sky130_fd_sc_hd__a22o_1 _2993_ (.A1(\weights_inst.data_out[3] ),
    .A2(_0654_),
    .B1(_0658_),
    .B2(\fsm_inst.done ),
    .X(net44));
 sky130_fd_sc_hd__and2_1 _2994_ (.A(\weights_inst.data_out[4] ),
    .B(_0654_),
    .X(_0659_));
 sky130_fd_sc_hd__buf_1 _2995_ (.A(_0659_),
    .X(net45));
 sky130_fd_sc_hd__and2_1 _2996_ (.A(\weights_inst.data_out[5] ),
    .B(_0654_),
    .X(_0660_));
 sky130_fd_sc_hd__buf_1 _2997_ (.A(_0660_),
    .X(net46));
 sky130_fd_sc_hd__and2_1 _2998_ (.A(\weights_inst.data_out[6] ),
    .B(_0654_),
    .X(_0662_));
 sky130_fd_sc_hd__buf_1 _2999_ (.A(_0662_),
    .X(net47));
 sky130_fd_sc_hd__and2_1 _3000_ (.A(\weights_inst.data_out[7] ),
    .B(_0654_),
    .X(_0663_));
 sky130_fd_sc_hd__buf_1 _3001_ (.A(_0663_),
    .X(net48));
 sky130_fd_sc_hd__and2_1 _3002_ (.A(\weights_inst.data_out[8] ),
    .B(_0654_),
    .X(_0664_));
 sky130_fd_sc_hd__buf_1 _3003_ (.A(_0664_),
    .X(net49));
 sky130_fd_sc_hd__and2_1 _3004_ (.A(\weights_inst.data_out[9] ),
    .B(_0654_),
    .X(_0665_));
 sky130_fd_sc_hd__buf_1 _3005_ (.A(_0665_),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_2 _3006_ (.A(net55),
    .X(_0666_));
 sky130_fd_sc_hd__and2_1 _3007_ (.A(\weights_inst.data_out[10] ),
    .B(_0666_),
    .X(_0668_));
 sky130_fd_sc_hd__buf_1 _3008_ (.A(_0668_),
    .X(net21));
 sky130_fd_sc_hd__and2_1 _3009_ (.A(\weights_inst.data_out[11] ),
    .B(_0666_),
    .X(_0669_));
 sky130_fd_sc_hd__buf_1 _3010_ (.A(_0669_),
    .X(net22));
 sky130_fd_sc_hd__and2_1 _3011_ (.A(\weights_inst.data_out[12] ),
    .B(_0666_),
    .X(_0670_));
 sky130_fd_sc_hd__buf_1 _3012_ (.A(_0670_),
    .X(net23));
 sky130_fd_sc_hd__and2_1 _3013_ (.A(\weights_inst.data_out[13] ),
    .B(_0666_),
    .X(_0671_));
 sky130_fd_sc_hd__buf_1 _3014_ (.A(_0671_),
    .X(net24));
 sky130_fd_sc_hd__and2_1 _3015_ (.A(\weights_inst.data_out[14] ),
    .B(_0666_),
    .X(_0672_));
 sky130_fd_sc_hd__buf_1 _3016_ (.A(_0672_),
    .X(net25));
 sky130_fd_sc_hd__and2_1 _3017_ (.A(\weights_inst.data_out[15] ),
    .B(_0666_),
    .X(_0674_));
 sky130_fd_sc_hd__buf_1 _3018_ (.A(_0674_),
    .X(net26));
 sky130_fd_sc_hd__and2_1 _3019_ (.A(\weights_inst.data_out[16] ),
    .B(_0666_),
    .X(_0675_));
 sky130_fd_sc_hd__buf_1 _3020_ (.A(_0675_),
    .X(net27));
 sky130_fd_sc_hd__and2_1 _3021_ (.A(\weights_inst.data_out[17] ),
    .B(_0666_),
    .X(_0676_));
 sky130_fd_sc_hd__buf_1 _3022_ (.A(_0676_),
    .X(net28));
 sky130_fd_sc_hd__and2_1 _3023_ (.A(\weights_inst.data_out[18] ),
    .B(_0666_),
    .X(_0677_));
 sky130_fd_sc_hd__buf_1 _3024_ (.A(_0677_),
    .X(net29));
 sky130_fd_sc_hd__and2_1 _3025_ (.A(\weights_inst.data_out[19] ),
    .B(_0666_),
    .X(_0678_));
 sky130_fd_sc_hd__buf_1 _3026_ (.A(_0678_),
    .X(net30));
 sky130_fd_sc_hd__and2_1 _3027_ (.A(\weights_inst.data_out[20] ),
    .B(net55),
    .X(_0680_));
 sky130_fd_sc_hd__buf_1 _3028_ (.A(_0680_),
    .X(net32));
 sky130_fd_sc_hd__and2_1 _3029_ (.A(\weights_inst.data_out[21] ),
    .B(net55),
    .X(_0681_));
 sky130_fd_sc_hd__buf_1 _3030_ (.A(_0681_),
    .X(net33));
 sky130_fd_sc_hd__and2_1 _3031_ (.A(\weights_inst.data_out[22] ),
    .B(net55),
    .X(_0682_));
 sky130_fd_sc_hd__buf_1 _3032_ (.A(_0682_),
    .X(net34));
 sky130_fd_sc_hd__and2_1 _3033_ (.A(\weights_inst.data_out[23] ),
    .B(net55),
    .X(_0683_));
 sky130_fd_sc_hd__buf_2 _3034_ (.A(_0683_),
    .X(net43));
 sky130_fd_sc_hd__and3b_1 _3035_ (.A_N(\fsm_inst.current_state[1] ),
    .B(\fsm_inst.current_state[0] ),
    .C(\fsm_inst.current_state[2] ),
    .X(_0684_));
 sky130_fd_sc_hd__clkbuf_1 _3036_ (.A(_0684_),
    .X(_0000_));
 sky130_fd_sc_hd__and3b_1 _3037_ (.A_N(\fsm_inst.current_state[0] ),
    .B(\fsm_inst.current_state[2] ),
    .C(\fsm_inst.current_state[1] ),
    .X(_0686_));
 sky130_fd_sc_hd__clkbuf_1 _3038_ (.A(_0686_),
    .X(_0001_));
 sky130_fd_sc_hd__and3_1 _3039_ (.A(\fsm_inst.current_state[1] ),
    .B(\fsm_inst.current_state[0] ),
    .C(\fsm_inst.current_state[2] ),
    .X(_0687_));
 sky130_fd_sc_hd__clkbuf_1 _3040_ (.A(_0687_),
    .X(_0002_));
 sky130_fd_sc_hd__inv_2 _3041_ (.A(net13),
    .Y(_0688_));
 sky130_fd_sc_hd__a21oi_1 _3042_ (.A1(net13),
    .A2(net14),
    .B1(net15),
    .Y(_0689_));
 sky130_fd_sc_hd__nor3b_1 _3043_ (.A(net14),
    .B(net15),
    .C_N(net16),
    .Y(_0690_));
 sky130_fd_sc_hd__o21ba_1 _3044_ (.A1(net16),
    .A2(_0689_),
    .B1_N(_0690_),
    .X(_0691_));
 sky130_fd_sc_hd__inv_2 _3045_ (.A(net18),
    .Y(_0692_));
 sky130_fd_sc_hd__or3_1 _3046_ (.A(\fsm_inst.current_state[1] ),
    .B(\fsm_inst.current_state[0] ),
    .C(\fsm_inst.current_state[2] ),
    .X(_0693_));
 sky130_fd_sc_hd__or4_2 _3047_ (.A(_0692_),
    .B(_0420_),
    .C(_0657_),
    .D(_0693_),
    .X(_0695_));
 sky130_fd_sc_hd__and3b_1 _3048_ (.A_N(net16),
    .B(net15),
    .C(net14),
    .X(_0696_));
 sky130_fd_sc_hd__a31o_1 _3049_ (.A1(\fsm_inst.current_state[1] ),
    .A2(_0688_),
    .A3(_0696_),
    .B1(\fsm_inst.current_state[2] ),
    .X(_0697_));
 sky130_fd_sc_hd__a21bo_1 _3050_ (.A1(\fsm_inst.current_state[0] ),
    .A2(_0697_),
    .B1_N(_0693_),
    .X(_0698_));
 sky130_fd_sc_hd__o31ai_1 _3051_ (.A1(_0688_),
    .A2(_0691_),
    .A3(_0695_),
    .B1(_0698_),
    .Y(\fsm_inst.next_state[0] ));
 sky130_fd_sc_hd__xnor2_1 _3052_ (.A(\fsm_inst.current_state[1] ),
    .B(\fsm_inst.current_state[0] ),
    .Y(_0699_));
 sky130_fd_sc_hd__o31ai_1 _3053_ (.A1(net14),
    .A2(_0691_),
    .A3(_0695_),
    .B1(_0699_),
    .Y(\fsm_inst.next_state[1] ));
 sky130_fd_sc_hd__nor2_1 _3054_ (.A(_0696_),
    .B(_0690_),
    .Y(_0700_));
 sky130_fd_sc_hd__a21oi_1 _3055_ (.A1(net13),
    .A2(_0690_),
    .B1(\fsm_inst.current_state[0] ),
    .Y(_0701_));
 sky130_fd_sc_hd__a21oi_1 _3056_ (.A1(\fsm_inst.current_state[1] ),
    .A2(\fsm_inst.current_state[0] ),
    .B1(\fsm_inst.current_state[2] ),
    .Y(_0702_));
 sky130_fd_sc_hd__a211o_1 _3057_ (.A1(\fsm_inst.current_state[1] ),
    .A2(_0701_),
    .B1(_0702_),
    .C1(_0002_),
    .X(_0704_));
 sky130_fd_sc_hd__o21ai_1 _3058_ (.A1(_0695_),
    .A2(_0700_),
    .B1(_0704_),
    .Y(\fsm_inst.next_state[2] ));
 sky130_fd_sc_hd__buf_4 _3059_ (.A(net1),
    .X(_0705_));
 sky130_fd_sc_hd__inv_2 _3060_ (.A(_0705_),
    .Y(_0028_));
 sky130_fd_sc_hd__inv_2 _3061_ (.A(_0705_),
    .Y(_0029_));
 sky130_fd_sc_hd__inv_2 _3062_ (.A(_0705_),
    .Y(_0030_));
 sky130_fd_sc_hd__inv_2 _3063_ (.A(_0705_),
    .Y(_0031_));
 sky130_fd_sc_hd__inv_2 _3064_ (.A(_0705_),
    .Y(_0032_));
 sky130_fd_sc_hd__inv_2 _3065_ (.A(_0705_),
    .Y(_0033_));
 sky130_fd_sc_hd__inv_2 _3066_ (.A(_0705_),
    .Y(_0034_));
 sky130_fd_sc_hd__inv_2 _3067_ (.A(_0705_),
    .Y(_0035_));
 sky130_fd_sc_hd__inv_2 _3068_ (.A(_0705_),
    .Y(_0036_));
 sky130_fd_sc_hd__inv_2 _3069_ (.A(_0705_),
    .Y(_0037_));
 sky130_fd_sc_hd__buf_4 _3070_ (.A(net1),
    .X(_0707_));
 sky130_fd_sc_hd__inv_2 _3071_ (.A(_0707_),
    .Y(_0038_));
 sky130_fd_sc_hd__inv_2 _3072_ (.A(_0707_),
    .Y(_0039_));
 sky130_fd_sc_hd__inv_2 _3073_ (.A(_0707_),
    .Y(_0040_));
 sky130_fd_sc_hd__inv_2 _3074_ (.A(_0707_),
    .Y(_0041_));
 sky130_fd_sc_hd__inv_2 _3075_ (.A(_0707_),
    .Y(_0042_));
 sky130_fd_sc_hd__inv_2 _3076_ (.A(_0707_),
    .Y(_0043_));
 sky130_fd_sc_hd__inv_2 _3077_ (.A(_0707_),
    .Y(_0044_));
 sky130_fd_sc_hd__inv_2 _3078_ (.A(_0707_),
    .Y(_0045_));
 sky130_fd_sc_hd__inv_2 _3079_ (.A(_0707_),
    .Y(_0046_));
 sky130_fd_sc_hd__inv_2 _3080_ (.A(_0707_),
    .Y(_0047_));
 sky130_fd_sc_hd__buf_4 _3081_ (.A(net1),
    .X(_0709_));
 sky130_fd_sc_hd__inv_2 _3082_ (.A(_0709_),
    .Y(_0048_));
 sky130_fd_sc_hd__inv_2 _3083_ (.A(_0709_),
    .Y(_0049_));
 sky130_fd_sc_hd__inv_2 _3084_ (.A(_0709_),
    .Y(_0050_));
 sky130_fd_sc_hd__inv_2 _3085_ (.A(_0709_),
    .Y(_0051_));
 sky130_fd_sc_hd__inv_2 _3086_ (.A(_0709_),
    .Y(_0052_));
 sky130_fd_sc_hd__inv_2 _3087_ (.A(_0709_),
    .Y(_0053_));
 sky130_fd_sc_hd__inv_2 _3088_ (.A(_0709_),
    .Y(_0054_));
 sky130_fd_sc_hd__inv_2 _3089_ (.A(_0709_),
    .Y(_0055_));
 sky130_fd_sc_hd__inv_2 _3090_ (.A(_0709_),
    .Y(_0056_));
 sky130_fd_sc_hd__inv_2 _3091_ (.A(_0709_),
    .Y(_0057_));
 sky130_fd_sc_hd__inv_2 _3092_ (.A(net1),
    .Y(_0058_));
 sky130_fd_sc_hd__dfrtp_1 _3093_ (.CLK(clknet_2_1__leaf_wb_clk_i),
    .D(_0003_),
    .RESET_B(_0028_),
    .Q(net19));
 sky130_fd_sc_hd__dfrtp_1 _3094_ (.CLK(clknet_2_0__leaf_wb_clk_i),
    .D(_0001_),
    .RESET_B(_0029_),
    .Q(\fsm_inst.batch_norm_en ));
 sky130_fd_sc_hd__dfrtp_1 _3095_ (.CLK(clknet_2_1__leaf_wb_clk_i),
    .D(_0002_),
    .RESET_B(_0030_),
    .Q(\fsm_inst.done ));
 sky130_fd_sc_hd__dfrtp_1 _3096_ (.CLK(clknet_2_1__leaf_wb_clk_i),
    .D(_0000_),
    .RESET_B(_0031_),
    .Q(\fsm_inst.cnn_en ));
 sky130_fd_sc_hd__dfrtp_4 _3097_ (.CLK(clknet_2_1__leaf_wb_clk_i),
    .D(net61),
    .RESET_B(_0032_),
    .Q(\fsm_inst.current_state[0] ));
 sky130_fd_sc_hd__dfrtp_4 _3098_ (.CLK(clknet_2_1__leaf_wb_clk_i),
    .D(net63),
    .RESET_B(_0033_),
    .Q(\fsm_inst.current_state[1] ));
 sky130_fd_sc_hd__dfrtp_1 _3099_ (.CLK(clknet_2_1__leaf_wb_clk_i),
    .D(net86),
    .RESET_B(_0034_),
    .Q(\fsm_inst.current_state[2] ));
 sky130_fd_sc_hd__dfrtp_1 _3100_ (.CLK(clknet_2_0__leaf_wb_clk_i),
    .D(_0004_),
    .RESET_B(_0035_),
    .Q(\weights_inst.data_out[0] ));
 sky130_fd_sc_hd__dfrtp_1 _3101_ (.CLK(clknet_2_1__leaf_wb_clk_i),
    .D(_0015_),
    .RESET_B(_0036_),
    .Q(\weights_inst.data_out[1] ));
 sky130_fd_sc_hd__dfrtp_1 _3102_ (.CLK(clknet_2_0__leaf_wb_clk_i),
    .D(_0019_),
    .RESET_B(_0037_),
    .Q(\weights_inst.data_out[2] ));
 sky130_fd_sc_hd__dfrtp_1 _3103_ (.CLK(clknet_2_0__leaf_wb_clk_i),
    .D(_0021_),
    .RESET_B(_0038_),
    .Q(\weights_inst.data_out[3] ));
 sky130_fd_sc_hd__dfrtp_1 _3104_ (.CLK(clknet_2_0__leaf_wb_clk_i),
    .D(_0022_),
    .RESET_B(_0039_),
    .Q(\weights_inst.data_out[4] ));
 sky130_fd_sc_hd__dfrtp_1 _3105_ (.CLK(clknet_2_3__leaf_wb_clk_i),
    .D(_0023_),
    .RESET_B(_0040_),
    .Q(\weights_inst.data_out[5] ));
 sky130_fd_sc_hd__dfrtp_1 _3106_ (.CLK(clknet_2_2__leaf_wb_clk_i),
    .D(_0024_),
    .RESET_B(_0041_),
    .Q(\weights_inst.data_out[6] ));
 sky130_fd_sc_hd__dfrtp_1 _3107_ (.CLK(clknet_2_0__leaf_wb_clk_i),
    .D(_0025_),
    .RESET_B(_0042_),
    .Q(\weights_inst.data_out[7] ));
 sky130_fd_sc_hd__dfrtp_1 _3108_ (.CLK(clknet_2_3__leaf_wb_clk_i),
    .D(_0026_),
    .RESET_B(_0043_),
    .Q(\weights_inst.data_out[8] ));
 sky130_fd_sc_hd__dfrtp_1 _3109_ (.CLK(clknet_2_2__leaf_wb_clk_i),
    .D(_0027_),
    .RESET_B(_0044_),
    .Q(\weights_inst.data_out[9] ));
 sky130_fd_sc_hd__dfrtp_1 _3110_ (.CLK(clknet_2_2__leaf_wb_clk_i),
    .D(_0005_),
    .RESET_B(_0045_),
    .Q(\weights_inst.data_out[10] ));
 sky130_fd_sc_hd__dfrtp_1 _3111_ (.CLK(clknet_2_2__leaf_wb_clk_i),
    .D(_0006_),
    .RESET_B(_0046_),
    .Q(\weights_inst.data_out[11] ));
 sky130_fd_sc_hd__dfrtp_1 _3112_ (.CLK(clknet_2_3__leaf_wb_clk_i),
    .D(_0007_),
    .RESET_B(_0047_),
    .Q(\weights_inst.data_out[12] ));
 sky130_fd_sc_hd__dfrtp_1 _3113_ (.CLK(clknet_2_2__leaf_wb_clk_i),
    .D(_0008_),
    .RESET_B(_0048_),
    .Q(\weights_inst.data_out[13] ));
 sky130_fd_sc_hd__dfrtp_1 _3114_ (.CLK(clknet_2_3__leaf_wb_clk_i),
    .D(_0009_),
    .RESET_B(_0049_),
    .Q(\weights_inst.data_out[14] ));
 sky130_fd_sc_hd__dfrtp_1 _3115_ (.CLK(clknet_2_2__leaf_wb_clk_i),
    .D(_0010_),
    .RESET_B(_0050_),
    .Q(\weights_inst.data_out[15] ));
 sky130_fd_sc_hd__dfrtp_1 _3116_ (.CLK(clknet_2_3__leaf_wb_clk_i),
    .D(_0011_),
    .RESET_B(_0051_),
    .Q(\weights_inst.data_out[16] ));
 sky130_fd_sc_hd__dfrtp_1 _3117_ (.CLK(clknet_2_2__leaf_wb_clk_i),
    .D(_0012_),
    .RESET_B(_0052_),
    .Q(\weights_inst.data_out[17] ));
 sky130_fd_sc_hd__dfrtp_1 _3118_ (.CLK(clknet_2_3__leaf_wb_clk_i),
    .D(_0013_),
    .RESET_B(_0053_),
    .Q(\weights_inst.data_out[18] ));
 sky130_fd_sc_hd__dfrtp_1 _3119_ (.CLK(clknet_2_3__leaf_wb_clk_i),
    .D(_0014_),
    .RESET_B(_0054_),
    .Q(\weights_inst.data_out[19] ));
 sky130_fd_sc_hd__dfrtp_1 _3120_ (.CLK(clknet_2_2__leaf_wb_clk_i),
    .D(_0016_),
    .RESET_B(_0055_),
    .Q(\weights_inst.data_out[20] ));
 sky130_fd_sc_hd__dfrtp_1 _3121_ (.CLK(clknet_2_3__leaf_wb_clk_i),
    .D(_0017_),
    .RESET_B(_0056_),
    .Q(\weights_inst.data_out[21] ));
 sky130_fd_sc_hd__dfrtp_1 _3122_ (.CLK(clknet_2_2__leaf_wb_clk_i),
    .D(_0018_),
    .RESET_B(_0057_),
    .Q(\weights_inst.data_out[22] ));
 sky130_fd_sc_hd__dfrtp_1 _3123_ (.CLK(clknet_2_3__leaf_wb_clk_i),
    .D(_0020_),
    .RESET_B(_0058_),
    .Q(\weights_inst.data_out[23] ));
 sky130_fd_sc_hd__buf_1 _3125_ (.A(net43),
    .X(net35));
 sky130_fd_sc_hd__buf_1 _3126_ (.A(net43),
    .X(net36));
 sky130_fd_sc_hd__buf_1 _3127_ (.A(net43),
    .X(net37));
 sky130_fd_sc_hd__buf_1 _3128_ (.A(net43),
    .X(net38));
 sky130_fd_sc_hd__buf_1 _3129_ (.A(net43),
    .X(net39));
 sky130_fd_sc_hd__buf_1 _3130_ (.A(net43),
    .X(net40));
 sky130_fd_sc_hd__buf_1 _3131_ (.A(net43),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_wb_clk_i (.A(wb_clk_i),
    .X(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(wbs_dat_i[0]),
    .X(net60));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(_0847_),
    .X(net69));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(_0862_),
    .X(net70));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(_0453_),
    .X(net71));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(_0454_),
    .X(net72));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(wbs_adr_i[1]),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_2 hold15 (.A(_0998_),
    .X(net74));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(_1074_),
    .X(net75));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(_1076_),
    .X(net76));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(wbs_adr_i[6]),
    .X(net77));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(_0846_),
    .X(net78));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\fsm_inst.next_state[0] ),
    .X(net61));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(wbs_adr_i[0]),
    .X(net79));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(wbs_adr_i[4]),
    .X(net80));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(wbs_adr_i[2]),
    .X(net81));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(wbs_adr_i[5]),
    .X(net82));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(wbs_adr_i[3]),
    .X(net83));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(wbs_adr_i[9]),
    .X(net84));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(net11),
    .X(net85));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\fsm_inst.next_state[2] ),
    .X(net86));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(net19),
    .X(net87));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(wbs_dat_i[1]),
    .X(net62));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\fsm_inst.next_state[1] ),
    .X(net63));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(wbs_adr_i[8]),
    .X(net64));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(net10),
    .X(net65));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold7 (.A(_0858_),
    .X(net66));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(_1157_),
    .X(net67));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(wbs_adr_i[7]),
    .X(net68));
 sky130_fd_sc_hd__buf_2 input1 (.A(wb_rst_i),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(net64),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(net84),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(wbs_cyc_i),
    .X(net12));
 sky130_fd_sc_hd__buf_1 input13 (.A(net60),
    .X(net13));
 sky130_fd_sc_hd__buf_1 input14 (.A(net62),
    .X(net14));
 sky130_fd_sc_hd__buf_1 input15 (.A(wbs_dat_i[2]),
    .X(net15));
 sky130_fd_sc_hd__buf_1 input16 (.A(wbs_dat_i[3]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(wbs_stb_i),
    .X(net17));
 sky130_fd_sc_hd__buf_1 input18 (.A(wbs_we_i),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(net79),
    .X(net2));
 sky130_fd_sc_hd__buf_4 input3 (.A(net73),
    .X(net3));
 sky130_fd_sc_hd__buf_4 input4 (.A(net81),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_2 input5 (.A(net83),
    .X(net5));
 sky130_fd_sc_hd__buf_4 input6 (.A(net80),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_4 input7 (.A(net82),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_2 input8 (.A(net77),
    .X(net8));
 sky130_fd_sc_hd__buf_4 input9 (.A(net68),
    .X(net9));
 sky130_fd_sc_hd__conb_1 kws_wrapper_59 (.LO(net59));
 sky130_fd_sc_hd__clkbuf_1 max_cap1 (.A(_0653_),
    .X(net88));
 sky130_fd_sc_hd__buf_2 max_cap51 (.A(_1422_),
    .X(net51));
 sky130_fd_sc_hd__buf_1 max_cap53 (.A(_0658_),
    .X(net53));
 sky130_fd_sc_hd__buf_4 max_cap54 (.A(_0880_),
    .X(net54));
 sky130_fd_sc_hd__buf_4 max_cap56 (.A(_0946_),
    .X(net56));
 sky130_fd_sc_hd__buf_4 max_cap57 (.A(_0766_),
    .X(net57));
 sky130_fd_sc_hd__buf_4 max_cap58 (.A(_0452_),
    .X(net58));
 sky130_fd_sc_hd__buf_12 output19 (.A(net19),
    .X(wbs_ack_o));
 sky130_fd_sc_hd__buf_12 output20 (.A(net20),
    .X(wbs_dat_o[0]));
 sky130_fd_sc_hd__buf_12 output21 (.A(net21),
    .X(wbs_dat_o[10]));
 sky130_fd_sc_hd__buf_12 output22 (.A(net22),
    .X(wbs_dat_o[11]));
 sky130_fd_sc_hd__buf_12 output23 (.A(net23),
    .X(wbs_dat_o[12]));
 sky130_fd_sc_hd__buf_12 output24 (.A(net24),
    .X(wbs_dat_o[13]));
 sky130_fd_sc_hd__buf_12 output25 (.A(net25),
    .X(wbs_dat_o[14]));
 sky130_fd_sc_hd__buf_12 output26 (.A(net26),
    .X(wbs_dat_o[15]));
 sky130_fd_sc_hd__buf_12 output27 (.A(net27),
    .X(wbs_dat_o[16]));
 sky130_fd_sc_hd__buf_12 output28 (.A(net28),
    .X(wbs_dat_o[17]));
 sky130_fd_sc_hd__buf_12 output29 (.A(net29),
    .X(wbs_dat_o[18]));
 sky130_fd_sc_hd__buf_12 output30 (.A(net30),
    .X(wbs_dat_o[19]));
 sky130_fd_sc_hd__buf_12 output31 (.A(net31),
    .X(wbs_dat_o[1]));
 sky130_fd_sc_hd__buf_12 output32 (.A(net32),
    .X(wbs_dat_o[20]));
 sky130_fd_sc_hd__buf_12 output33 (.A(net33),
    .X(wbs_dat_o[21]));
 sky130_fd_sc_hd__buf_12 output34 (.A(net34),
    .X(wbs_dat_o[22]));
 sky130_fd_sc_hd__buf_12 output35 (.A(net35),
    .X(wbs_dat_o[23]));
 sky130_fd_sc_hd__buf_12 output36 (.A(net36),
    .X(wbs_dat_o[24]));
 sky130_fd_sc_hd__buf_12 output37 (.A(net37),
    .X(wbs_dat_o[25]));
 sky130_fd_sc_hd__buf_12 output38 (.A(net38),
    .X(wbs_dat_o[26]));
 sky130_fd_sc_hd__buf_12 output39 (.A(net39),
    .X(wbs_dat_o[27]));
 sky130_fd_sc_hd__buf_12 output40 (.A(net40),
    .X(wbs_dat_o[28]));
 sky130_fd_sc_hd__buf_12 output41 (.A(net41),
    .X(wbs_dat_o[29]));
 sky130_fd_sc_hd__buf_12 output42 (.A(net42),
    .X(wbs_dat_o[2]));
 sky130_fd_sc_hd__buf_12 output43 (.A(net43),
    .X(wbs_dat_o[30]));
 sky130_fd_sc_hd__buf_12 output44 (.A(net44),
    .X(wbs_dat_o[3]));
 sky130_fd_sc_hd__buf_12 output45 (.A(net45),
    .X(wbs_dat_o[4]));
 sky130_fd_sc_hd__buf_12 output46 (.A(net46),
    .X(wbs_dat_o[5]));
 sky130_fd_sc_hd__buf_12 output47 (.A(net47),
    .X(wbs_dat_o[6]));
 sky130_fd_sc_hd__buf_12 output48 (.A(net48),
    .X(wbs_dat_o[7]));
 sky130_fd_sc_hd__buf_12 output49 (.A(net49),
    .X(wbs_dat_o[8]));
 sky130_fd_sc_hd__buf_12 output50 (.A(net50),
    .X(wbs_dat_o[9]));
 sky130_fd_sc_hd__buf_4 wire52 (.A(_0773_),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_2 wire55 (.A(net88),
    .X(net55));
 assign wbs_dat_o[31] = net59;
endmodule

