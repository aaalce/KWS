* NGSPICE file created from kws_wrapper.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_4 abstract view
.subckt sky130_fd_sc_hd__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_4 abstract view
.subckt sky130_fd_sc_hd__and2b_4 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_1 abstract view
.subckt sky130_fd_sc_hd__o311ai_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_4 abstract view
.subckt sky130_fd_sc_hd__a311o_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_4 abstract view
.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

.subckt kws_wrapper VGND VPWR wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10]
+ wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16]
+ wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21]
+ wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27]
+ wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3]
+ wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i
+ wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14]
+ wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1]
+ wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25]
+ wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30]
+ wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8]
+ wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13]
+ wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19]
+ wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24]
+ wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2]
+ wbs_dat_o[30] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8]
+ wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
+ wbs_dat_o[31]
XFILLER_0_94_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3086_ _0709_ VGND VGND VPWR VPWR _0052_ sky130_fd_sc_hd__inv_2
X_2106_ _0763_ _0891_ VGND VGND VPWR VPWR _1247_ sky130_fd_sc_hd__and2_4
XFILLER_0_89_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2037_ _0811_ _1172_ _1174_ _1177_ _1178_ VGND VGND VPWR VPWR _1179_ sky130_fd_sc_hd__o311a_1
XFILLER_0_76_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2939_ _0838_ _0599_ _0600_ _0604_ _0841_ VGND VGND VPWR VPWR _0605_ sky130_fd_sc_hd__a311o_2
XFILLER_0_45_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2724_ _0911_ _0974_ _1094_ VGND VGND VPWR VPWR _0378_ sky130_fd_sc_hd__or3_1
XFILLER_0_42_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2655_ _0843_ _0308_ _0310_ VGND VGND VPWR VPWR _0311_ sky130_fd_sc_hd__or3_1
X_1606_ _0750_ VGND VGND VPWR VPWR _0751_ sky130_fd_sc_hd__buf_4
X_2586_ _1109_ _0925_ _1354_ _0243_ _0978_ VGND VGND VPWR VPWR _0244_ sky130_fd_sc_hd__o311a_1
X_1537_ net7 net5 VGND VGND VPWR VPWR _0462_ sky130_fd_sc_hd__and2_1
XTAP_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3069_ _0705_ VGND VGND VPWR VPWR _0037_ sky130_fd_sc_hd__inv_2
XFILLER_0_92_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2440_ _1274_ _0733_ _1130_ _0100_ _1198_ VGND VGND VPWR VPWR _0101_ sky130_fd_sc_hd__o311a_1
XFILLER_0_51_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2371_ _0957_ _1283_ _1448_ _1507_ _0963_ VGND VGND VPWR VPWR _1508_ sky130_fd_sc_hd__o311a_1
XFILLER_0_75_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2707_ _0791_ _1358_ _0922_ VGND VGND VPWR VPWR _0362_ sky130_fd_sc_hd__a21o_1
XFILLER_0_71_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2638_ _0878_ _0973_ _0130_ _0922_ VGND VGND VPWR VPWR _0295_ sky130_fd_sc_hd__a211o_1
X_2569_ _0917_ _1066_ _0942_ VGND VGND VPWR VPWR _0227_ sky130_fd_sc_hd__a21o_1
XFILLER_0_100_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_364 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1940_ _0799_ VGND VGND VPWR VPWR _1083_ sky130_fd_sc_hd__buf_4
XFILLER_0_16_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1871_ _0784_ VGND VGND VPWR VPWR _1015_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_28_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2423_ _1443_ _0080_ VGND VGND VPWR VPWR _0085_ sky130_fd_sc_hd__and2b_1
XFILLER_0_20_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2354_ _0728_ _0829_ VGND VGND VPWR VPWR _1491_ sky130_fd_sc_hd__nor2_4
X_2285_ _1000_ _1229_ _1176_ _1140_ VGND VGND VPWR VPWR _1424_ sky130_fd_sc_hd__a211o_1
XFILLER_0_79_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2070_ _0824_ _0815_ _1097_ _1199_ _1211_ VGND VGND VPWR VPWR _1212_ sky130_fd_sc_hd__a221o_1
XFILLER_0_88_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2972_ _1291_ _0639_ _0608_ VGND VGND VPWR VPWR _0640_ sky130_fd_sc_hd__o21ai_1
XTAP_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1923_ _0757_ _0720_ _1007_ VGND VGND VPWR VPWR _1067_ sky130_fd_sc_hd__or3_4
XFILLER_0_8_339 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1854_ _0717_ net3 VGND VGND VPWR VPWR _0998_ sky130_fd_sc_hd__xor2_1
XFILLER_0_4_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1785_ _0742_ _0830_ VGND VGND VPWR VPWR _0930_ sky130_fd_sc_hd__nor2_4
XFILLER_0_97_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2406_ _1110_ _0886_ _0879_ _1365_ VGND VGND VPWR VPWR _0068_ sky130_fd_sc_hd__o211a_1
X_2337_ _0728_ _1391_ VGND VGND VPWR VPWR _1475_ sky130_fd_sc_hd__nor2_4
XFILLER_0_34_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2268_ _0718_ _0763_ _0732_ VGND VGND VPWR VPWR _1407_ sky130_fd_sc_hd__and3_4
X_2199_ _0800_ _0890_ _1118_ VGND VGND VPWR VPWR _1339_ sky130_fd_sc_hd__or3_1
XFILLER_0_67_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1570_ net58 _0714_ VGND VGND VPWR VPWR _0715_ sky130_fd_sc_hd__xor2_4
XANTENNA_5 _0215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2122_ _0791_ _1044_ _1262_ VGND VGND VPWR VPWR _1263_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_83_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2053_ _1164_ _1171_ _1179_ _1194_ VGND VGND VPWR VPWR _1195_ sky130_fd_sc_hd__o31a_1
XFILLER_0_88_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2955_ _0621_ VGND VGND VPWR VPWR _0018_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2886_ _0786_ _0868_ _1202_ _1140_ VGND VGND VPWR VPWR _0547_ sky130_fd_sc_hd__a211o_1
XFILLER_0_44_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1906_ _1003_ _1015_ VGND VGND VPWR VPWR _1050_ sky130_fd_sc_hd__nor2_4
XFILLER_0_72_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1837_ _0944_ _0979_ _0980_ VGND VGND VPWR VPWR _0981_ sky130_fd_sc_hd__or3_1
X_1768_ _0881_ _0829_ _0785_ VGND VGND VPWR VPWR _0913_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_12_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1699_ _0783_ _0792_ _0809_ _0840_ _0843_ VGND VGND VPWR VPWR _0844_ sky130_fd_sc_hd__a311o_1
XFILLER_0_40_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput42 net42 VGND VGND VPWR VPWR wbs_dat_o[2] sky130_fd_sc_hd__buf_12
Xoutput20 net20 VGND VGND VPWR VPWR wbs_dat_o[0] sky130_fd_sc_hd__buf_12
Xoutput31 net31 VGND VGND VPWR VPWR wbs_dat_o[1] sky130_fd_sc_hd__buf_12
XFILLER_0_101_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2740_ _1299_ _1323_ _0393_ _0752_ _1308_ VGND VGND VPWR VPWR _0394_ sky130_fd_sc_hd__o221a_1
XFILLER_0_81_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2671_ _1311_ _1097_ _1127_ _0824_ _1264_ VGND VGND VPWR VPWR _0327_ sky130_fd_sc_hd__a221o_1
XFILLER_0_54_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1622_ _0765_ net57 VGND VGND VPWR VPWR _0767_ sky130_fd_sc_hd__nor2_8
XFILLER_0_10_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1553_ _0602_ _0623_ VGND VGND VPWR VPWR _0634_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_22_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3085_ _0709_ VGND VGND VPWR VPWR _0051_ sky130_fd_sc_hd__inv_2
X_2105_ _1233_ _1245_ VGND VGND VPWR VPWR _1246_ sky130_fd_sc_hd__nor2_2
XFILLER_0_89_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2036_ _0914_ VGND VGND VPWR VPWR _1178_ sky130_fd_sc_hd__buf_4
XFILLER_0_49_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_423 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2938_ _0601_ _0603_ _0776_ VGND VGND VPWR VPWR _0604_ sky130_fd_sc_hd__o21a_1
XFILLER_0_17_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2869_ _1343_ _0996_ _0940_ _1261_ _1329_ VGND VGND VPWR VPWR _0530_ sky130_fd_sc_hd__o221ai_2
XFILLER_0_60_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_392 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2723_ _1347_ _0903_ _0919_ VGND VGND VPWR VPWR _0377_ sky130_fd_sc_hd__o21a_1
XFILLER_0_81_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2654_ _0816_ _1500_ _0309_ _1274_ _1178_ VGND VGND VPWR VPWR _0310_ sky130_fd_sc_hd__o221a_1
X_2585_ _1013_ _1206_ _0180_ _1011_ _0800_ VGND VGND VPWR VPWR _0243_ sky130_fd_sc_hd__a221o_1
XFILLER_0_22_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1605_ _0749_ VGND VGND VPWR VPWR _0750_ sky130_fd_sc_hd__buf_4
XFILLER_0_10_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1536_ net7 net5 VGND VGND VPWR VPWR _0452_ sky130_fd_sc_hd__xor2_4
XFILLER_0_89_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3068_ _0705_ VGND VGND VPWR VPWR _0036_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2019_ _1036_ VGND VGND VPWR VPWR _1161_ sky130_fd_sc_hd__buf_4
XFILLER_0_92_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2370_ _0916_ _0815_ _1506_ _0970_ _1028_ VGND VGND VPWR VPWR _1507_ sky130_fd_sc_hd__a221o_1
XFILLER_0_75_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_170 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2706_ _0999_ _0815_ _1183_ _1028_ VGND VGND VPWR VPWR _0361_ sky130_fd_sc_hd__a211o_1
X_2637_ _0292_ _0293_ _0957_ VGND VGND VPWR VPWR _0294_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2568_ _0824_ _0815_ _1475_ _1211_ VGND VGND VPWR VPWR _0226_ sky130_fd_sc_hd__a211o_1
XFILLER_0_10_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2499_ _0810_ _1050_ _1077_ VGND VGND VPWR VPWR _0159_ sky130_fd_sc_hd__or3_1
XFILLER_0_97_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1870_ _1012_ _1013_ VGND VGND VPWR VPWR _1014_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2422_ _0074_ _0083_ _1161_ VGND VGND VPWR VPWR _0084_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_19_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2353_ _1078_ _1059_ VGND VGND VPWR VPWR _1490_ sky130_fd_sc_hd__nor2_1
X_2284_ _0452_ _0813_ net51 _1232_ _1165_ VGND VGND VPWR VPWR _1423_ sky130_fd_sc_hd__a221o_1
XFILLER_0_79_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1999_ _1123_ _1001_ VGND VGND VPWR VPWR _1142_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_170 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2971_ _0824_ _0807_ _0130_ VGND VGND VPWR VPWR _0639_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_56_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1922_ _0784_ _0767_ VGND VGND VPWR VPWR _1066_ sky130_fd_sc_hd__nor2_4
XFILLER_0_16_107 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1853_ _0758_ _0996_ VGND VGND VPWR VPWR _0997_ sky130_fd_sc_hd__nor2_2
XFILLER_0_4_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1784_ _0851_ VGND VGND VPWR VPWR _0929_ sky130_fd_sc_hd__buf_4
XFILLER_0_24_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2405_ _0062_ _0066_ _1365_ VGND VGND VPWR VPWR _0067_ sky130_fd_sc_hd__a21oi_2
X_2336_ _0797_ _1084_ _1150_ _0835_ VGND VGND VPWR VPWR _1474_ sky130_fd_sc_hd__a211o_1
X_2267_ _1244_ _1181_ _1405_ _1310_ VGND VGND VPWR VPWR _1406_ sky130_fd_sc_hd__o211a_1
XFILLER_0_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2198_ _1042_ _1337_ _0935_ VGND VGND VPWR VPWR _1338_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_75_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold20 wbs_adr_i[0] VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_85_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_6 _0253_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2121_ _1261_ _0938_ VGND VGND VPWR VPWR _1262_ sky130_fd_sc_hd__nor2_1
XFILLER_0_83_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2052_ _0703_ _1186_ _1192_ _1193_ VGND VGND VPWR VPWR _1194_ sky130_fd_sc_hd__a211o_1
XFILLER_0_88_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2954_ _0859_ _0620_ VGND VGND VPWR VPWR _0621_ sky130_fd_sc_hd__and2_1
XFILLER_0_29_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2885_ _0970_ _1213_ _0744_ _0739_ VGND VGND VPWR VPWR _0546_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_17_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1905_ _0864_ VGND VGND VPWR VPWR _1049_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_4_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1836_ _0756_ _0820_ VGND VGND VPWR VPWR _0980_ sky130_fd_sc_hd__nor2_2
X_1767_ _0745_ _0732_ _0831_ VGND VGND VPWR VPWR _0912_ sky130_fd_sc_hd__and3_2
XFILLER_0_40_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1698_ _0842_ VGND VGND VPWR VPWR _0843_ sky130_fd_sc_hd__buf_4
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2319_ _0852_ _0727_ _0996_ VGND VGND VPWR VPWR _1457_ sky130_fd_sc_hd__and3_2
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput21 net21 VGND VGND VPWR VPWR wbs_dat_o[10] sky130_fd_sc_hd__buf_12
Xoutput32 net32 VGND VGND VPWR VPWR wbs_dat_o[20] sky130_fd_sc_hd__buf_12
Xoutput43 net43 VGND VGND VPWR VPWR wbs_dat_o[30] sky130_fd_sc_hd__buf_12
XFILLER_0_53_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2670_ _1345_ _0960_ _1059_ _0325_ _1287_ VGND VGND VPWR VPWR _0326_ sky130_fd_sc_hd__o311a_1
XFILLER_0_81_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1621_ _0717_ _0708_ VGND VGND VPWR VPWR _0766_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_41_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1552_ net9 _0613_ VGND VGND VPWR VPWR _0623_ sky130_fd_sc_hd__xnor2_4
X_2104_ _1123_ _0971_ _0970_ VGND VGND VPWR VPWR _1245_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_89_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3084_ _0709_ VGND VGND VPWR VPWR _0050_ sky130_fd_sc_hd__inv_2
X_2035_ _1049_ _1175_ _1176_ VGND VGND VPWR VPWR _1177_ sky130_fd_sc_hd__or3_1
XFILLER_0_89_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_360 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2937_ _0791_ _0805_ _1392_ _1078_ _0833_ VGND VGND VPWR VPWR _0603_ sky130_fd_sc_hd__o221a_1
XFILLER_0_94_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2868_ _0221_ _0528_ _1356_ VGND VGND VPWR VPWR _0529_ sky130_fd_sc_hd__o21a_1
XFILLER_0_60_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2799_ net72 VGND VGND VPWR VPWR _0013_ sky130_fd_sc_hd__buf_1
X_1819_ _0685_ VGND VGND VPWR VPWR _0963_ sky130_fd_sc_hd__buf_4
XFILLER_0_60_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2722_ _1158_ _0351_ _0352_ _0376_ _0859_ VGND VGND VPWR VPWR _0011_ sky130_fd_sc_hd__o311a_1
XFILLER_0_54_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2653_ _1016_ _1301_ VGND VGND VPWR VPWR _0309_ sky130_fd_sc_hd__nor2_1
X_2584_ _1298_ _0234_ _0235_ _0241_ VGND VGND VPWR VPWR _0242_ sky130_fd_sc_hd__o31ai_2
X_1604_ _0723_ VGND VGND VPWR VPWR _0749_ sky130_fd_sc_hd__clkbuf_4
X_1535_ net7 net9 VGND VGND VPWR VPWR _0441_ sky130_fd_sc_hd__xor2_4
XFILLER_0_10_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3067_ _0705_ VGND VGND VPWR VPWR _0035_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2018_ _0975_ _1159_ VGND VGND VPWR VPWR _1160_ sky130_fd_sc_hd__nand2_4
XFILLER_0_54_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2705_ _0273_ _0358_ _0359_ _1264_ VGND VGND VPWR VPWR _0360_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_42_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2636_ _1247_ _0289_ VGND VGND VPWR VPWR _0293_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2567_ _1256_ _0931_ _0146_ _0224_ _1193_ VGND VGND VPWR VPWR _0225_ sky130_fd_sc_hd__o311a_1
XFILLER_0_57_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2498_ _0852_ _1011_ _1025_ _0985_ VGND VGND VPWR VPWR _0158_ sky130_fd_sc_hd__a31o_1
XFILLER_0_97_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3119_ clknet_2_3__leaf_wb_clk_i _0014_ _0054_ VGND VGND VPWR VPWR weights_inst.data_out\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_300 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_388 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2421_ _0842_ _0078_ _0082_ VGND VGND VPWR VPWR _0083_ sky130_fd_sc_hd__or3b_2
X_2352_ _0816_ _0817_ _1448_ _1264_ VGND VGND VPWR VPWR _1489_ sky130_fd_sc_hd__a211o_1
XFILLER_0_19_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2283_ _0728_ _0720_ _1007_ VGND VGND VPWR VPWR _1422_ sky130_fd_sc_hd__nor3_4
XFILLER_0_19_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_439 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1998_ _0852_ _1041_ VGND VGND VPWR VPWR _1141_ sky130_fd_sc_hd__nor2_2
XFILLER_0_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2619_ _1198_ _0274_ _0275_ _0907_ VGND VGND VPWR VPWR _0276_ sky130_fd_sc_hd__a31o_1
XFILLER_0_65_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2970_ _0605_ _0637_ _1396_ VGND VGND VPWR VPWR _0638_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_29_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1921_ _0926_ _1064_ VGND VGND VPWR VPWR _1065_ sky130_fd_sc_hd__nand2_8
XFILLER_0_71_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1852_ _0718_ _0711_ VGND VGND VPWR VPWR _0996_ sky130_fd_sc_hd__nand2_8
XFILLER_0_4_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1783_ _0926_ _0802_ _0927_ VGND VGND VPWR VPWR _0928_ sky130_fd_sc_hd__and3_2
XFILLER_0_40_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2404_ _0706_ _0063_ _0064_ _0065_ _1164_ VGND VGND VPWR VPWR _0066_ sky130_fd_sc_hd__a311o_1
X_2335_ _0694_ _1471_ _1472_ VGND VGND VPWR VPWR _1473_ sky130_fd_sc_hd__and3_1
X_2266_ _1232_ _1311_ _0787_ _0801_ VGND VGND VPWR VPWR _1405_ sky130_fd_sc_hd__a211o_1
X_2197_ _1291_ _0722_ VGND VGND VPWR VPWR _1337_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold10 _0847_ VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 wbs_adr_i[4] VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_7 _0298_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2120_ _1083_ VGND VGND VPWR VPWR _1261_ sky130_fd_sc_hd__buf_4
X_2051_ _0841_ VGND VGND VPWR VPWR _1193_ sky130_fd_sc_hd__buf_4
XFILLER_0_88_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2953_ _0576_ _0589_ _0606_ _0619_ _1036_ _0848_ VGND VGND VPWR VPWR _0620_ sky130_fd_sc_hd__mux4_1
XFILLER_0_57_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1904_ _1040_ _0774_ _1042_ _1046_ _1047_ VGND VGND VPWR VPWR _1048_ sky130_fd_sc_hd__o311a_1
XFILLER_0_57_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2884_ _1193_ _0536_ _0539_ _0544_ _0860_ VGND VGND VPWR VPWR _0545_ sky130_fd_sc_hd__o311a_1
XFILLER_0_72_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1835_ _0918_ _0870_ VGND VGND VPWR VPWR _0979_ sky130_fd_sc_hd__nor2_1
X_1766_ _0910_ VGND VGND VPWR VPWR _0911_ sky130_fd_sc_hd__buf_4
XFILLER_0_12_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1697_ _0841_ VGND VGND VPWR VPWR _0842_ sky130_fd_sc_hd__buf_4
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2318_ _0743_ _1001_ VGND VGND VPWR VPWR _1456_ sky130_fd_sc_hd__nor2_1
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2249_ _1244_ _1326_ _1323_ _1387_ _1356_ VGND VGND VPWR VPWR _1388_ sky130_fd_sc_hd__o311a_1
XFILLER_0_95_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_450 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput22 net22 VGND VGND VPWR VPWR wbs_dat_o[11] sky130_fd_sc_hd__buf_12
Xoutput33 net33 VGND VGND VPWR VPWR wbs_dat_o[21] sky130_fd_sc_hd__buf_12
XFILLER_0_9_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput44 net44 VGND VGND VPWR VPWR wbs_dat_o[3] sky130_fd_sc_hd__buf_12
XFILLER_0_98_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_328 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_383 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1620_ _0731_ VGND VGND VPWR VPWR _0765_ sky130_fd_sc_hd__clkbuf_16
X_1551_ _0537_ _0570_ _0527_ VGND VGND VPWR VPWR _0613_ sky130_fd_sc_hd__a21boi_4
X_2103_ _1040_ VGND VGND VPWR VPWR _1244_ sky130_fd_sc_hd__buf_4
X_3083_ _0709_ VGND VGND VPWR VPWR _0049_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2034_ _0452_ _0947_ VGND VGND VPWR VPWR _1176_ sky130_fd_sc_hd__nor2_1
XFILLER_0_89_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2936_ _0745_ _1073_ _0257_ _0723_ VGND VGND VPWR VPWR _0601_ sky130_fd_sc_hd__o211a_1
XFILLER_0_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2867_ _0940_ _1487_ _0873_ VGND VGND VPWR VPWR _0528_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1818_ _0877_ _0961_ VGND VGND VPWR VPWR _0962_ sky130_fd_sc_hd__and2_1
X_2798_ net66 _0437_ net71 VGND VGND VPWR VPWR _0454_ sky130_fd_sc_hd__and3_1
X_1749_ _0806_ _0867_ _0893_ _0754_ VGND VGND VPWR VPWR _0894_ sky130_fd_sc_hd__a211o_1
XFILLER_0_40_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2721_ _0365_ _0375_ _1197_ VGND VGND VPWR VPWR _0376_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_81_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2652_ _1256_ _1475_ net52 _0307_ _0703_ VGND VGND VPWR VPWR _0308_ sky130_fd_sc_hd__o311a_1
XFILLER_0_22_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1603_ _0739_ _0744_ _0747_ VGND VGND VPWR VPWR _0748_ sky130_fd_sc_hd__a21o_1
X_2583_ _1310_ _0236_ _0238_ _0240_ _1318_ VGND VGND VPWR VPWR _0241_ sky130_fd_sc_hd__a311o_1
X_1534_ net87 _0420_ VGND VGND VPWR VPWR _0003_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_51 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3066_ _0705_ VGND VGND VPWR VPWR _0034_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2017_ _0741_ _0812_ VGND VGND VPWR VPWR _1159_ sky130_fd_sc_hd__nor2_2
XFILLER_0_18_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2919_ _1099_ _1407_ _0749_ VGND VGND VPWR VPWR _0583_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_18_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_364 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2704_ _0880_ _1016_ _1073_ _1077_ VGND VGND VPWR VPWR _0359_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2635_ _0970_ _1506_ _1324_ _0929_ VGND VGND VPWR VPWR _0292_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2566_ _0755_ _0966_ _1305_ VGND VGND VPWR VPWR _0224_ sky130_fd_sc_hd__or3_1
XFILLER_0_49_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2497_ _1198_ _0152_ _0153_ _0156_ VGND VGND VPWR VPWR _0157_ sky130_fd_sc_hd__a31o_1
X_3118_ clknet_2_3__leaf_wb_clk_i _0013_ _0053_ VGND VGND VPWR VPWR weights_inst.data_out\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3049_ fsm_inst.current_state\[1\] _0688_ _0696_ fsm_inst.current_state\[2\] VGND
+ VGND VPWR VPWR _0697_ sky130_fd_sc_hd__a31o_1
XFILLER_0_81_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_312 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2420_ _0810_ _1160_ _0079_ _0081_ _0838_ VGND VGND VPWR VPWR _0082_ sky130_fd_sc_hd__a311o_1
XFILLER_0_86_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2351_ _0810_ _1050_ _1410_ _1487_ VGND VGND VPWR VPWR _1488_ sky130_fd_sc_hd__or4_1
X_2282_ _0739_ _0744_ _0816_ _1078_ _0923_ VGND VGND VPWR VPWR _1421_ sky130_fd_sc_hd__a221o_1
XFILLER_0_79_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1997_ _0984_ VGND VGND VPWR VPWR _1140_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_15_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2618_ _1060_ _1030_ _0997_ _1314_ VGND VGND VPWR VPWR _0275_ sky130_fd_sc_hd__or4_1
XFILLER_0_11_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2549_ _1348_ _0733_ _1524_ _0207_ _1310_ VGND VGND VPWR VPWR _0208_ sky130_fd_sc_hd__o311a_1
XFILLER_0_97_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1920_ _0735_ _0999_ VGND VGND VPWR VPWR _1064_ sky130_fd_sc_hd__nor2_8
XFILLER_0_84_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1851_ _0952_ _0969_ _0982_ _0994_ _0860_ VGND VGND VPWR VPWR _0995_ sky130_fd_sc_hd__o311a_1
XFILLER_0_71_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1782_ _0742_ _0886_ VGND VGND VPWR VPWR _0927_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2403_ _1225_ _1294_ _1253_ _1400_ _1178_ VGND VGND VPWR VPWR _0065_ sky130_fd_sc_hd__o221a_1
X_2334_ _0828_ _1084_ _1127_ _0823_ _0864_ VGND VGND VPWR VPWR _1472_ sky130_fd_sc_hd__a221o_1
X_2265_ _0889_ _1400_ _1402_ _1403_ _0935_ VGND VGND VPWR VPWR _1404_ sky130_fd_sc_hd__o221a_1
X_2196_ _1182_ _1334_ _1335_ VGND VGND VPWR VPWR _1336_ sky130_fd_sc_hd__o21a_1
XFILLER_0_79_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_61 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold11 _0862_ VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__dlygate4sd3_1
Xhold22 wbs_adr_i[2] VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_8 _0340_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2050_ _1187_ _1189_ _1191_ _0875_ _0914_ VGND VGND VPWR VPWR _1192_ sky130_fd_sc_hd__o221a_1
XFILLER_0_76_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2952_ _1193_ _0609_ _0611_ _0618_ VGND VGND VPWR VPWR _0619_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_29_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1903_ _0838_ VGND VGND VPWR VPWR _1047_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_72_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2883_ _0661_ _0541_ _0543_ VGND VGND VPWR VPWR _0544_ sky130_fd_sc_hd__or3_1
X_1834_ _0777_ VGND VGND VPWR VPWR _0978_ sky130_fd_sc_hd__buf_4
XFILLER_0_4_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1765_ _0834_ VGND VGND VPWR VPWR _0910_ sky130_fd_sc_hd__buf_4
XFILLER_0_40_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1696_ _0516_ _0580_ VGND VGND VPWR VPWR _0841_ sky130_fd_sc_hd__xnor2_4
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2317_ _0800_ _1001_ _1453_ _1454_ VGND VGND VPWR VPWR _1455_ sky130_fd_sc_hd__a31o_1
XFILLER_0_57_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2248_ _1229_ _0965_ _1230_ _0923_ VGND VGND VPWR VPWR _1387_ sky130_fd_sc_hd__a211o_1
XFILLER_0_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2179_ _1298_ _1304_ _1309_ _1319_ _1039_ VGND VGND VPWR VPWR _1320_ sky130_fd_sc_hd__o311a_1
XFILLER_0_73_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput34 net34 VGND VGND VPWR VPWR wbs_dat_o[22] sky130_fd_sc_hd__buf_12
Xoutput23 net23 VGND VGND VPWR VPWR wbs_dat_o[12] sky130_fd_sc_hd__buf_12
Xoutput45 net45 VGND VGND VPWR VPWR wbs_dat_o[4] sky130_fd_sc_hd__buf_12
XFILLER_0_98_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_395 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1550_ _0591_ VGND VGND VPWR VPWR _0602_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2102_ _1193_ VGND VGND VPWR VPWR _1243_ sky130_fd_sc_hd__buf_4
XFILLER_0_27_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3082_ _0709_ VGND VGND VPWR VPWR _0048_ sky130_fd_sc_hd__inv_2
X_2033_ _0877_ _1173_ VGND VGND VPWR VPWR _1175_ sky130_fd_sc_hd__nor2_4
XFILLER_0_72_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2935_ _0771_ _0389_ _0956_ VGND VGND VPWR VPWR _0600_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_57_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2866_ _0522_ _0525_ _0673_ VGND VGND VPWR VPWR _0526_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_32_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1817_ _0771_ _0959_ VGND VGND VPWR VPWR _0961_ sky130_fd_sc_hd__nand2_4
X_2797_ _0449_ _0451_ _0863_ VGND VGND VPWR VPWR _0453_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1748_ _0758_ _0892_ VGND VGND VPWR VPWR _0893_ sky130_fd_sc_hd__nor2_2
X_1679_ _0823_ VGND VGND VPWR VPWR _0824_ sky130_fd_sc_hd__buf_4
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2720_ _1039_ _0367_ _0369_ _0374_ _1243_ VGND VGND VPWR VPWR _0375_ sky130_fd_sc_hd__o311a_1
XFILLER_0_14_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2651_ _1083_ _1009_ _0266_ VGND VGND VPWR VPWR _0307_ sky130_fd_sc_hd__or3_1
XFILLER_0_54_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1602_ _0741_ _0745_ _0746_ VGND VGND VPWR VPWR _0747_ sky130_fd_sc_hd__and3_2
XFILLER_0_22_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2582_ _0957_ _1326_ _1501_ _0239_ _0778_ VGND VGND VPWR VPWR _0240_ sky130_fd_sc_hd__o311a_1
X_1533_ net17 net12 VGND VGND VPWR VPWR _0420_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3065_ _0705_ VGND VGND VPWR VPWR _0033_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2016_ _0849_ VGND VGND VPWR VPWR _1158_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_49_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2918_ _0579_ _0581_ _0694_ VGND VGND VPWR VPWR _0582_ sky130_fd_sc_hd__a21o_1
XFILLER_0_33_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2849_ _0911_ _0827_ _1359_ VGND VGND VPWR VPWR _0508_ sky130_fd_sc_hd__or3b_1
XFILLER_0_60_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2703_ _0834_ _0899_ VGND VGND VPWR VPWR _0358_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2634_ _1348_ _1079_ _0289_ _0290_ _1310_ VGND VGND VPWR VPWR _0291_ sky130_fd_sc_hd__o311a_1
XFILLER_0_2_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2565_ _0811_ _1470_ _0221_ _0222_ _0907_ VGND VGND VPWR VPWR _0223_ sky130_fd_sc_hd__o311a_1
XFILLER_0_10_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2496_ _1235_ _1066_ _1166_ _0155_ _0950_ VGND VGND VPWR VPWR _0156_ sky130_fd_sc_hd__o311a_1
X_3117_ clknet_2_2__leaf_wb_clk_i _0012_ _0052_ VGND VGND VPWR VPWR weights_inst.data_out\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_3048_ net16 net15 net14 VGND VGND VPWR VPWR _0696_ sky130_fd_sc_hd__and3b_1
XFILLER_0_65_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_143 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2350_ _0825_ _0820_ _1025_ VGND VGND VPWR VPWR _1487_ sky130_fd_sc_hd__and3_1
XFILLER_0_19_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2281_ _1281_ _1247_ _1417_ _1419_ _1356_ VGND VGND VPWR VPWR _1420_ sky130_fd_sc_hd__o311a_1
XFILLER_0_87_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1996_ _1091_ _1135_ _1138_ VGND VGND VPWR VPWR _1139_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_27_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2617_ _1232_ _0786_ _0867_ _0273_ _0873_ VGND VGND VPWR VPWR _0274_ sky130_fd_sc_hd__a311o_1
XFILLER_0_11_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2548_ _1049_ _0733_ _1183_ _1265_ VGND VGND VPWR VPWR _0207_ sky130_fd_sc_hd__or4_1
X_2479_ _1264_ _1111_ _1500_ _0138_ VGND VGND VPWR VPWR _0139_ sky130_fd_sc_hd__o31a_1
XFILLER_0_97_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1850_ _0978_ _0986_ _0987_ _0992_ _0993_ VGND VGND VPWR VPWR _0994_ sky130_fd_sc_hd__a311o_1
XFILLER_0_21_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1781_ _0757_ VGND VGND VPWR VPWR _0926_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_52_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2402_ _1256_ _0980_ _1283_ VGND VGND VPWR VPWR _0064_ sky130_fd_sc_hd__or3_1
X_2333_ _1013_ _1205_ _1470_ _0754_ VGND VGND VPWR VPWR _1471_ sky130_fd_sc_hd__a211o_1
X_2264_ _1180_ VGND VGND VPWR VPWR _1403_ sky130_fd_sc_hd__buf_4
XFILLER_0_79_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2195_ _1211_ VGND VGND VPWR VPWR _1335_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_216 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1979_ _0751_ _1118_ _1119_ _0978_ _1121_ VGND VGND VPWR VPWR _1122_ sky130_fd_sc_hd__o311a_1
XFILLER_0_43_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold12 _0453_ VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 wbs_adr_i[5] VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_9 _0374_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2951_ _0778_ _0612_ _0614_ _0617_ VGND VGND VPWR VPWR _0618_ sky130_fd_sc_hd__a31o_1
XFILLER_0_84_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1902_ _1019_ _1043_ _0916_ _1045_ _0800_ VGND VGND VPWR VPWR _1046_ sky130_fd_sc_hd__a221o_1
XFILLER_0_72_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2882_ _1187_ _0542_ _0694_ VGND VGND VPWR VPWR _0543_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_72_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1833_ _0975_ _0971_ _0976_ VGND VGND VPWR VPWR _0977_ sky130_fd_sc_hd__and3_2
X_1764_ _0863_ _0908_ VGND VGND VPWR VPWR _0909_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1695_ _0811_ _0822_ _0837_ _0839_ VGND VGND VPWR VPWR _0840_ sky130_fd_sc_hd__o211a_4
XFILLER_0_0_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2316_ _0787_ _1188_ _0869_ _1236_ _0984_ VGND VGND VPWR VPWR _1454_ sky130_fd_sc_hd__o221a_1
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2247_ _1250_ _1385_ VGND VGND VPWR VPWR _1386_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2178_ _1310_ _1312_ _1313_ _1317_ _1318_ VGND VGND VPWR VPWR _1319_ sky130_fd_sc_hd__a311o_1
XFILLER_0_95_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput24 net24 VGND VGND VPWR VPWR wbs_dat_o[13] sky130_fd_sc_hd__buf_12
XFILLER_0_31_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput46 net46 VGND VGND VPWR VPWR wbs_dat_o[5] sky130_fd_sc_hd__buf_12
Xoutput35 net35 VGND VGND VPWR VPWR wbs_dat_o[23] sky130_fd_sc_hd__buf_12
XFILLER_0_98_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2101_ _1158_ _1196_ _1241_ _1242_ VGND VGND VPWR VPWR _0021_ sky130_fd_sc_hd__o211a_1
X_3081_ net1 VGND VGND VPWR VPWR _0709_ sky130_fd_sc_hd__buf_4
X_2032_ _1117_ _1173_ VGND VGND VPWR VPWR _1174_ sky130_fd_sc_hd__nor2_2
XFILLER_0_77_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2934_ _1127_ _1422_ _0910_ _1232_ VGND VGND VPWR VPWR _0599_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_72_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2865_ _1278_ _0523_ _0524_ VGND VGND VPWR VPWR _0525_ sky130_fd_sc_hd__and3_2
XFILLER_0_72_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1816_ _0745_ _0790_ _0959_ VGND VGND VPWR VPWR _0960_ sky130_fd_sc_hd__and3_2
X_2796_ _0787_ _0901_ _0450_ _0860_ VGND VGND VPWR VPWR _0451_ sky130_fd_sc_hd__o31a_1
X_1747_ _0891_ VGND VGND VPWR VPWR _0892_ sky130_fd_sc_hd__buf_4
X_1678_ _0719_ VGND VGND VPWR VPWR _0823_ sky130_fd_sc_hd__buf_4
XFILLER_0_68_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_311 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2650_ _0706_ _0301_ _0302_ _0305_ _1164_ VGND VGND VPWR VPWR _0306_ sky130_fd_sc_hd__a311o_1
XFILLER_0_42_506 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1601_ _0718_ _0731_ VGND VGND VPWR VPWR _0746_ sky130_fd_sc_hd__nand2_2
X_2581_ _0803_ _1072_ _0146_ _0985_ VGND VGND VPWR VPWR _0239_ sky130_fd_sc_hd__a211o_1
XFILLER_0_10_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3064_ _0705_ VGND VGND VPWR VPWR _0032_ sky130_fd_sc_hd__inv_2
X_2015_ net67 VGND VGND VPWR VPWR _0019_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2917_ _0928_ _0450_ _0800_ VGND VGND VPWR VPWR _0581_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_45_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2848_ _0706_ _0502_ _0506_ VGND VGND VPWR VPWR _0507_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_5_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2779_ _0749_ _0898_ _1457_ VGND VGND VPWR VPWR _0433_ sky130_fd_sc_hd__or3_1
XFILLER_0_41_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2702_ _1281_ _1300_ _0214_ _0356_ _1285_ VGND VGND VPWR VPWR _0357_ sky130_fd_sc_hd__o311a_1
XFILLER_0_27_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2633_ _1347_ _1097_ _1259_ VGND VGND VPWR VPWR _0290_ sky130_fd_sc_hd__a21o_1
XFILLER_0_2_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2564_ _0824_ _0827_ _1099_ _0803_ _1235_ VGND VGND VPWR VPWR _0222_ sky130_fd_sc_hd__a221o_1
XFILLER_0_100_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2495_ _0806_ _1399_ _0154_ _0956_ VGND VGND VPWR VPWR _0155_ sky130_fd_sc_hd__a211o_1
XFILLER_0_65_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3116_ clknet_2_3__leaf_wb_clk_i _0011_ _0051_ VGND VGND VPWR VPWR weights_inst.data_out\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_3047_ _0692_ _0420_ _0657_ _0693_ VGND VGND VPWR VPWR _0695_ sky130_fd_sc_hd__or4_2
XFILLER_0_65_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_196 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2280_ _1078_ _1229_ _1418_ _0801_ VGND VGND VPWR VPWR _1419_ sky130_fd_sc_hd__a211o_1
XFILLER_0_99_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1995_ _1136_ _0788_ _1137_ _1028_ VGND VGND VPWR VPWR _1138_ sky130_fd_sc_hd__a211o_1
XFILLER_0_15_369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2616_ _1136_ _1213_ VGND VGND VPWR VPWR _0273_ sky130_fd_sc_hd__nor2_2
XFILLER_0_23_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2547_ _1273_ _0197_ _0199_ _0205_ _1396_ VGND VGND VPWR VPWR _0206_ sky130_fd_sc_hd__o311a_1
XFILLER_0_11_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2478_ _0956_ _1094_ _0137_ VGND VGND VPWR VPWR _0138_ sky130_fd_sc_hd__or3_1
XFILLER_0_76_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1780_ _0825_ _0728_ _0924_ VGND VGND VPWR VPWR _0925_ sky130_fd_sc_hd__and3_4
XFILLER_0_97_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2401_ _1276_ _0811_ _1085_ VGND VGND VPWR VPWR _0063_ sky130_fd_sc_hd__or3b_2
X_2332_ _0740_ _0854_ _0897_ VGND VGND VPWR VPWR _1470_ sky130_fd_sc_hd__and3_2
X_2263_ _1189_ _1401_ VGND VGND VPWR VPWR _1402_ sky130_fd_sc_hd__and2b_1
X_2194_ _0763_ _0891_ _0927_ VGND VGND VPWR VPWR _1334_ sky130_fd_sc_hd__and3_2
XFILLER_0_46_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1978_ _1120_ _0739_ _0836_ VGND VGND VPWR VPWR _1121_ sky130_fd_sc_hd__a21o_1
XFILLER_0_43_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold13 _0454_ VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 wbs_adr_i[3] VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_214 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2950_ _0685_ _0615_ _0616_ _0661_ VGND VGND VPWR VPWR _0617_ sky130_fd_sc_hd__a31o_2
XFILLER_0_32_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2881_ _0767_ _0931_ _1028_ VGND VGND VPWR VPWR _0542_ sky130_fd_sc_hd__o21ai_1
X_1901_ _1015_ _1044_ VGND VGND VPWR VPWR _1045_ sky130_fd_sc_hd__nor2_2
X_1832_ _0742_ net57 VGND VGND VPWR VPWR _0976_ sky130_fd_sc_hd__nand2_8
XFILLER_0_25_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1763_ _0874_ _0884_ _0895_ _0906_ _0782_ _0907_ VGND VGND VPWR VPWR _0908_ sky130_fd_sc_hd__mux4_1
XFILLER_0_25_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1694_ _0838_ VGND VGND VPWR VPWR _0839_ sky130_fd_sc_hd__buf_4
XFILLER_0_40_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2315_ _0721_ _0829_ VGND VGND VPWR VPWR _1453_ sky130_fd_sc_hd__nand2_1
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2246_ _0811_ _0966_ _1172_ _1384_ VGND VGND VPWR VPWR _1385_ sky130_fd_sc_hd__o31a_1
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2177_ _0993_ VGND VGND VPWR VPWR _1318_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_18_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput25 net25 VGND VGND VPWR VPWR wbs_dat_o[14] sky130_fd_sc_hd__buf_12
XFILLER_0_31_467 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput36 net36 VGND VGND VPWR VPWR wbs_dat_o[24] sky130_fd_sc_hd__buf_12
Xoutput47 net47 VGND VGND VPWR VPWR wbs_dat_o[6] sky130_fd_sc_hd__buf_12
XFILLER_0_3_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2100_ net66 VGND VGND VPWR VPWR _1242_ sky130_fd_sc_hd__buf_2
X_3080_ _0707_ VGND VGND VPWR VPWR _0047_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2031_ _0772_ _0765_ _0741_ VGND VGND VPWR VPWR _1173_ sky130_fd_sc_hd__a21o_4
XFILLER_0_43_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2933_ _0593_ _0597_ VGND VGND VPWR VPWR _0598_ sky130_fd_sc_hd__nor2_1
XFILLER_0_72_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2864_ _0803_ _1099_ _1142_ _1040_ VGND VGND VPWR VPWR _0524_ sky130_fd_sc_hd__a211o_1
XFILLER_0_72_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1815_ _0958_ VGND VGND VPWR VPWR _0959_ sky130_fd_sc_hd__buf_4
XFILLER_0_32_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2795_ _0881_ _0797_ _0769_ VGND VGND VPWR VPWR _0450_ sky130_fd_sc_hd__a21oi_4
X_1746_ _0717_ _0708_ _0710_ VGND VGND VPWR VPWR _0891_ sky130_fd_sc_hd__or3_2
XFILLER_0_40_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1677_ _0816_ _0817_ _0821_ VGND VGND VPWR VPWR _0822_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_7_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2229_ _1183_ _1299_ _1366_ _1368_ _1308_ VGND VGND VPWR VPWR _1369_ sky130_fd_sc_hd__o311a_1
XFILLER_0_82_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1600_ _0727_ VGND VGND VPWR VPWR _0745_ sky130_fd_sc_hd__buf_4
XFILLER_0_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2580_ _0237_ _1379_ _1335_ VGND VGND VPWR VPWR _0238_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_10_448 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3063_ _0705_ VGND VGND VPWR VPWR _0031_ sky130_fd_sc_hd__inv_2
X_2014_ net66 _1108_ _1156_ VGND VGND VPWR VPWR _1157_ sky130_fd_sc_hd__and3_1
XFILLER_0_54_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2916_ _0855_ _0331_ _0985_ VGND VGND VPWR VPWR _0579_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_72_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_420 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2847_ _0783_ _0503_ _0504_ _1318_ VGND VGND VPWR VPWR _0506_ sky130_fd_sc_hd__a31o_1
XFILLER_0_60_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2778_ _1124_ _1491_ _1524_ _0922_ VGND VGND VPWR VPWR _0432_ sky130_fd_sc_hd__a211o_1
XFILLER_0_13_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1729_ _0760_ _0865_ _0867_ _0872_ _0873_ VGND VGND VPWR VPWR _0874_ sky130_fd_sc_hd__o32a_1
XFILLER_0_41_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_194 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2701_ _1367_ _0973_ _1410_ _0801_ VGND VGND VPWR VPWR _0356_ sky130_fd_sc_hd__a211o_1
XFILLER_0_15_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2632_ _0820_ _0924_ _0947_ VGND VGND VPWR VPWR _0289_ sky130_fd_sc_hd__and3_1
XFILLER_0_23_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2563_ _0770_ _1019_ _0983_ VGND VGND VPWR VPWR _0221_ sky130_fd_sc_hd__and3_2
XFILLER_0_2_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2494_ _0756_ _0745_ _0719_ VGND VGND VPWR VPWR _0154_ sky130_fd_sc_hd__and3_4
XFILLER_0_10_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3115_ clknet_2_2__leaf_wb_clk_i _0010_ _0050_ VGND VGND VPWR VPWR weights_inst.data_out\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_3046_ fsm_inst.current_state\[1\] fsm_inst.current_state\[0\] fsm_inst.current_state\[2\]
+ VGND VGND VPWR VPWR _0693_ sky130_fd_sc_hd__or3_1
XFILLER_0_77_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1994_ _0716_ _0738_ _0796_ VGND VGND VPWR VPWR _1137_ sky130_fd_sc_hd__and3_2
XFILLER_0_70_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2615_ _1281_ _0974_ _1443_ _0271_ VGND VGND VPWR VPWR _0272_ sky130_fd_sc_hd__o31a_1
XFILLER_0_30_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2546_ _0779_ _0200_ _0201_ _0204_ _0667_ VGND VGND VPWR VPWR _0205_ sky130_fd_sc_hd__a311o_1
X_2477_ _0757_ _0712_ _0965_ VGND VGND VPWR VPWR _0137_ sky130_fd_sc_hd__and3_4
XFILLER_0_48_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3029_ weights_inst.data_out\[21\] net55 VGND VGND VPWR VPWR _0681_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2400_ _1250_ _1531_ _0059_ _0061_ _1273_ VGND VGND VPWR VPWR _0062_ sky130_fd_sc_hd__a311o_1
XFILLER_0_24_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2331_ _0922_ _1466_ _1467_ _1468_ _0914_ VGND VGND VPWR VPWR _1469_ sky130_fd_sc_hd__o311a_1
X_2262_ _0802_ _1105_ VGND VGND VPWR VPWR _1401_ sky130_fd_sc_hd__nand2_1
X_2193_ _1328_ _1164_ _1332_ VGND VGND VPWR VPWR _1333_ sky130_fd_sc_hd__and3b_1
XFILLER_0_79_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1977_ _0975_ _1013_ VGND VGND VPWR VPWR _1120_ sky130_fd_sc_hd__nand2_2
XFILLER_0_55_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2529_ _1403_ _0919_ _1098_ _1278_ VGND VGND VPWR VPWR _0188_ sky130_fd_sc_hd__a31o_1
Xhold14 wbs_adr_i[1] VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 wbs_adr_i[9] VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1900_ _0828_ _0868_ VGND VGND VPWR VPWR _1044_ sky130_fd_sc_hd__nor2_4
X_2880_ _0964_ _1026_ _1168_ _0540_ _0838_ VGND VGND VPWR VPWR _0541_ sky130_fd_sc_hd__o311a_1
XTAP_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1831_ _0939_ VGND VGND VPWR VPWR _0975_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_25_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1762_ _0661_ VGND VGND VPWR VPWR _0907_ sky130_fd_sc_hd__buf_4
XFILLER_0_25_476 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1693_ _0685_ VGND VGND VPWR VPWR _0838_ sky130_fd_sc_hd__buf_4
XFILLER_0_0_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2314_ _0934_ _1450_ _1451_ _0841_ VGND VGND VPWR VPWR _1452_ sky130_fd_sc_hd__a31o_1
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2245_ _1049_ _1050_ _1350_ VGND VGND VPWR VPWR _1384_ sky130_fd_sc_hd__or3b_1
XFILLER_0_57_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2176_ _0957_ _1103_ _1255_ _1316_ _0778_ VGND VGND VPWR VPWR _1317_ sky130_fd_sc_hd__o311a_1
XFILLER_0_79_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput26 net26 VGND VGND VPWR VPWR wbs_dat_o[15] sky130_fd_sc_hd__buf_12
Xoutput37 net37 VGND VGND VPWR VPWR wbs_dat_o[25] sky130_fd_sc_hd__buf_12
Xoutput48 net48 VGND VGND VPWR VPWR wbs_dat_o[7] sky130_fd_sc_hd__buf_12
XFILLER_0_101_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2030_ _0877_ _1159_ VGND VGND VPWR VPWR _1172_ sky130_fd_sc_hd__nor2_2
XFILLER_0_69_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2932_ _0595_ _0596_ _0914_ VGND VGND VPWR VPWR _0597_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_57_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2863_ _1467_ _0875_ _1160_ VGND VGND VPWR VPWR _0523_ sky130_fd_sc_hd__or3b_1
XFILLER_0_72_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1814_ net2 net3 VGND VGND VPWR VPWR _0958_ sky130_fd_sc_hd__or2_1
X_2794_ _0667_ _0439_ _0442_ _0448_ _1036_ VGND VGND VPWR VPWR _0449_ sky130_fd_sc_hd__o311a_2
X_1745_ _0784_ _0746_ VGND VGND VPWR VPWR _0890_ sky130_fd_sc_hd__nor2_8
XFILLER_0_7_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1676_ _0713_ _0819_ _0820_ VGND VGND VPWR VPWR _0821_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_68_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2228_ _1019_ _1072_ _0965_ _1367_ _0751_ VGND VGND VPWR VPWR _1368_ sky130_fd_sc_hd__a221o_1
XFILLER_0_95_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2159_ _0878_ _0961_ VGND VGND VPWR VPWR _1300_ sky130_fd_sc_hd__nor2_2
XFILLER_0_95_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3131_ net43 VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__buf_1
XFILLER_0_38_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3062_ _0705_ VGND VGND VPWR VPWR _0030_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2013_ _1134_ _1155_ _0849_ VGND VGND VPWR VPWR _1156_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_54_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2915_ _1235_ _1141_ _1500_ _0577_ _0694_ VGND VGND VPWR VPWR _0578_ sky130_fd_sc_hd__o311ai_4
XFILLER_0_72_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2846_ _1232_ _1127_ _1410_ _1261_ VGND VGND VPWR VPWR _0504_ sky130_fd_sc_hd__a211o_1
XFILLER_0_5_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2777_ _0983_ _0948_ _1112_ _1140_ VGND VGND VPWR VPWR _0431_ sky130_fd_sc_hd__a211o_1
XFILLER_0_13_243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1728_ _0754_ VGND VGND VPWR VPWR _0873_ sky130_fd_sc_hd__buf_4
XFILLER_0_41_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1659_ _0718_ _0711_ VGND VGND VPWR VPWR _0804_ sky130_fd_sc_hd__nor2_1
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2700_ _1410_ _0353_ _0354_ VGND VGND VPWR VPWR _0355_ sky130_fd_sc_hd__o21a_1
X_2631_ _1345_ _0798_ _1512_ _0287_ _0935_ VGND VGND VPWR VPWR _0288_ sky130_fd_sc_hd__o311a_1
XFILLER_0_23_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2562_ _0860_ _0803_ _1020_ VGND VGND VPWR VPWR _0220_ sky130_fd_sc_hd__and3_1
XFILLER_0_23_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2493_ _1060_ _1050_ _1190_ _1410_ VGND VGND VPWR VPWR _0153_ sky130_fd_sc_hd__or4_1
XFILLER_0_4_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3114_ clknet_2_3__leaf_wb_clk_i _0009_ _0049_ VGND VGND VPWR VPWR weights_inst.data_out\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_3045_ net18 VGND VGND VPWR VPWR _0692_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2829_ _1053_ _1073_ _1165_ _0827_ VGND VGND VPWR VPWR _0487_ sky130_fd_sc_hd__a211o_1
XFILLER_0_5_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_382 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1993_ _1015_ VGND VGND VPWR VPWR _1136_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_70_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2614_ _1366_ _0270_ _1345_ VGND VGND VPWR VPWR _0271_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_42_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2545_ _0202_ _0203_ _1115_ VGND VGND VPWR VPWR _0204_ sky130_fd_sc_hd__o21a_2
XFILLER_0_76_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2476_ _1036_ _0737_ _1343_ VGND VGND VPWR VPWR _0136_ sky130_fd_sc_hd__or3_1
XFILLER_0_76_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3028_ _0680_ VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__buf_1
XFILLER_0_93_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_168 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2330_ _0834_ _0888_ _1301_ VGND VGND VPWR VPWR _1468_ sky130_fd_sc_hd__or3_1
X_2261_ _1011_ _1399_ VGND VGND VPWR VPWR _1400_ sky130_fd_sc_hd__nor2_1
X_2192_ _0789_ _0876_ _1329_ _1331_ _0915_ VGND VGND VPWR VPWR _1332_ sky130_fd_sc_hd__a221o_1
XFILLER_0_46_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1976_ _0918_ _0817_ VGND VGND VPWR VPWR _1119_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2528_ _1345_ _1344_ _0186_ VGND VGND VPWR VPWR _0187_ sky130_fd_sc_hd__and3_1
Xhold26 net11 VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__dlygate4sd3_1
X_2459_ _1273_ _0112_ _0114_ _0119_ _1161_ VGND VGND VPWR VPWR _0120_ sky130_fd_sc_hd__o311a_1
Xhold15 _0998_ VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_97_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_46 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1830_ _0970_ _0971_ _0973_ VGND VGND VPWR VPWR _0974_ sky130_fd_sc_hd__and3_2
XFILLER_0_13_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1761_ _0898_ _0900_ _0905_ VGND VGND VPWR VPWR _0906_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_25_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1692_ _0824_ _0827_ _0832_ _0836_ VGND VGND VPWR VPWR _0837_ sky130_fd_sc_hd__a211o_1
XFILLER_0_40_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2313_ _0835_ _1249_ _1085_ VGND VGND VPWR VPWR _1451_ sky130_fd_sc_hd__or3b_1
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2244_ _0817_ _1379_ _0913_ VGND VGND VPWR VPWR _1383_ sky130_fd_sc_hd__a21o_1
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2175_ _0824_ _1314_ _1315_ _0985_ VGND VGND VPWR VPWR _1316_ sky130_fd_sc_hd__a211o_1
XFILLER_0_79_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1959_ _1082_ _1087_ _1093_ _1101_ _0950_ _0842_ VGND VGND VPWR VPWR _1102_ sky130_fd_sc_hd__mux4_2
XFILLER_0_31_425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput49 net49 VGND VGND VPWR VPWR wbs_dat_o[8] sky130_fd_sc_hd__buf_12
Xoutput27 net27 VGND VGND VPWR VPWR wbs_dat_o[16] sky130_fd_sc_hd__buf_12
Xoutput38 net38 VGND VGND VPWR VPWR wbs_dat_o[26] sky130_fd_sc_hd__buf_12
XFILLER_0_98_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2931_ _1117_ _0896_ _0887_ _0864_ VGND VGND VPWR VPWR _0596_ sky130_fd_sc_hd__a211o_1
XFILLER_0_57_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2862_ _1345_ _0270_ _0303_ _0521_ _0779_ VGND VGND VPWR VPWR _0522_ sky130_fd_sc_hd__o311a_1
X_2793_ _0978_ _0443_ _0445_ _0447_ _0842_ VGND VGND VPWR VPWR _0448_ sky130_fd_sc_hd__a311o_1
XFILLER_0_53_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1813_ _0956_ VGND VGND VPWR VPWR _0957_ sky130_fd_sc_hd__buf_4
X_1744_ _0864_ _0888_ VGND VGND VPWR VPWR _0889_ sky130_fd_sc_hd__or2_2
XFILLER_0_4_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1675_ _0740_ VGND VGND VPWR VPWR _0820_ sky130_fd_sc_hd__buf_4
XFILLER_0_68_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2227_ _0975_ VGND VGND VPWR VPWR _1367_ sky130_fd_sc_hd__buf_4
XFILLER_0_84_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2158_ _0755_ _0882_ VGND VGND VPWR VPWR _1299_ sky130_fd_sc_hd__nand2_4
XFILLER_0_95_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2089_ _1229_ _1020_ _1230_ _0945_ VGND VGND VPWR VPWR _1231_ sky130_fd_sc_hd__a211o_1
XFILLER_0_48_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_366 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3130_ net43 VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__buf_1
X_3061_ _0705_ VGND VGND VPWR VPWR _0029_ sky130_fd_sc_hd__inv_2
X_2012_ _1039_ _1154_ VGND VGND VPWR VPWR _1155_ sky130_fd_sc_hd__nor2_1
XFILLER_0_77_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2914_ _1111_ _0209_ _1049_ VGND VGND VPWR VPWR _0577_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_72_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2845_ _0721_ _0739_ _1106_ _1165_ VGND VGND VPWR VPWR _0503_ sky130_fd_sc_hd__a211o_1
XFILLER_0_72_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2776_ _1264_ _1190_ _1202_ _0429_ _1047_ VGND VGND VPWR VPWR _0430_ sky130_fd_sc_hd__o311a_1
XFILLER_0_53_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1727_ _0868_ _0869_ _0871_ VGND VGND VPWR VPWR _0872_ sky130_fd_sc_hd__o21a_1
XFILLER_0_41_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1658_ _0802_ VGND VGND VPWR VPWR _0803_ sky130_fd_sc_hd__buf_8
XFILLER_0_95_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1589_ _0725_ _0733_ VGND VGND VPWR VPWR _0734_ sky130_fd_sc_hd__nor2_2
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_111 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2630_ _0983_ _1314_ _1335_ VGND VGND VPWR VPWR _0287_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_42_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2561_ _1158_ _0194_ _0219_ _1242_ VGND VGND VPWR VPWR _0007_ sky130_fd_sc_hd__o211a_1
XFILLER_0_23_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2492_ _1367_ _1113_ _0917_ _1467_ _0725_ VGND VGND VPWR VPWR _0152_ sky130_fd_sc_hd__a311o_1
XFILLER_0_23_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3113_ clknet_2_2__leaf_wb_clk_i _0008_ _0048_ VGND VGND VPWR VPWR weights_inst.data_out\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_3044_ net16 _0689_ _0690_ VGND VGND VPWR VPWR _0691_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_77_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2828_ _1347_ _1073_ VGND VGND VPWR VPWR _0486_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2759_ _0407_ _0412_ _1039_ VGND VGND VPWR VPWR _0413_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_41_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1992_ _0881_ _0786_ VGND VGND VPWR VPWR _1135_ sky130_fd_sc_hd__nor2_2
XFILLER_0_70_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_199 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2613_ _0770_ _1219_ _0976_ VGND VGND VPWR VPWR _0270_ sky130_fd_sc_hd__and3_1
XFILLER_0_30_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2544_ _0737_ _1011_ _0093_ _0922_ VGND VGND VPWR VPWR _0203_ sky130_fd_sc_hd__o211a_1
X_2475_ _1322_ _0121_ _0134_ _0135_ _0859_ VGND VGND VPWR VPWR _0005_ sky130_fd_sc_hd__o221a_1
XFILLER_0_76_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3027_ weights_inst.data_out\[20\] net55 VGND VGND VPWR VPWR _0680_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_420 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2260_ _0741_ _0996_ VGND VGND VPWR VPWR _1399_ sky130_fd_sc_hd__nand2_8
X_2191_ _1056_ _1330_ VGND VGND VPWR VPWR _1331_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1975_ _1117_ _0983_ VGND VGND VPWR VPWR _1118_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2527_ _0877_ _0887_ _0896_ VGND VGND VPWR VPWR _0186_ sky130_fd_sc_hd__or3_4
XFILLER_0_11_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2458_ _1278_ _0116_ _0118_ _0907_ VGND VGND VPWR VPWR _0119_ sky130_fd_sc_hd__a211o_1
Xhold16 _1074_ VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__dlygate4sd3_1
Xhold27 fsm_inst.next_state\[2\] VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__dlygate4sd3_1
X_2389_ _0957_ _1043_ _1523_ _1525_ _0978_ VGND VGND VPWR VPWR _1526_ sky130_fd_sc_hd__o311a_1
XFILLER_0_19_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_59 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1760_ _0869_ _0901_ _0902_ _0799_ _0904_ VGND VGND VPWR VPWR _0905_ sky130_fd_sc_hd__o221a_1
XFILLER_0_52_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1691_ _0835_ VGND VGND VPWR VPWR _0836_ sky130_fd_sc_hd__buf_4
XFILLER_0_52_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2312_ _1448_ _1449_ _1235_ VGND VGND VPWR VPWR _1450_ sky130_fd_sc_hd__o21ai_1
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2243_ _1322_ _1364_ _1382_ _1242_ VGND VGND VPWR VPWR _0023_ sky130_fd_sc_hd__o211a_1
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2174_ _1123_ _0819_ _1041_ VGND VGND VPWR VPWR _1315_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_94_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1958_ _1094_ _1096_ _1098_ _1100_ VGND VGND VPWR VPWR _1101_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_71_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1889_ _0756_ _1030_ _1032_ _0864_ VGND VGND VPWR VPWR _1033_ sky130_fd_sc_hd__a211o_1
XFILLER_0_31_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput28 net28 VGND VGND VPWR VPWR wbs_dat_o[17] sky130_fd_sc_hd__buf_12
Xoutput39 net39 VGND VGND VPWR VPWR wbs_dat_o[27] sky130_fd_sc_hd__buf_12
XFILLER_0_11_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2930_ _1432_ _0594_ _1028_ VGND VGND VPWR VPWR _0595_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_43_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2861_ _1400_ _0725_ _0722_ VGND VGND VPWR VPWR _0521_ sky130_fd_sc_hd__or3b_1
XFILLER_0_38_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1812_ _0749_ VGND VGND VPWR VPWR _0956_ sky130_fd_sc_hd__buf_4
X_2792_ _0944_ _0821_ _0146_ _0446_ _0838_ VGND VGND VPWR VPWR _0447_ sky130_fd_sc_hd__o311a_1
X_1743_ _0757_ _0887_ VGND VGND VPWR VPWR _0888_ sky130_fd_sc_hd__nor2_4
XFILLER_0_53_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1674_ _0818_ VGND VGND VPWR VPWR _0819_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2226_ _1064_ _1275_ VGND VGND VPWR VPWR _1366_ sky130_fd_sc_hd__nor2_1
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2157_ _1193_ VGND VGND VPWR VPWR _1298_ sky130_fd_sc_hd__buf_4
XFILLER_0_95_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2088_ _0926_ _0738_ _0924_ VGND VGND VPWR VPWR _1230_ sky130_fd_sc_hd__and3_2
XFILLER_0_48_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_223 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3060_ _0705_ VGND VGND VPWR VPWR _0028_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2011_ _1139_ _1145_ _1149_ _1153_ _0778_ _0907_ VGND VGND VPWR VPWR _1154_ sky130_fd_sc_hd__mux4_2
XFILLER_0_77_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2913_ _1125_ _0124_ VGND VGND VPWR VPWR _0576_ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2844_ _0828_ _1244_ _1084_ _0501_ VGND VGND VPWR VPWR _0502_ sky130_fd_sc_hd__a31o_1
XFILLER_0_72_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2775_ _0917_ _1152_ _1253_ VGND VGND VPWR VPWR _0429_ sky130_fd_sc_hd__a21o_1
X_1726_ _0768_ _0805_ _0870_ VGND VGND VPWR VPWR _0871_ sky130_fd_sc_hd__or3b_4
X_1657_ _0732_ VGND VGND VPWR VPWR _0802_ sky130_fd_sc_hd__buf_4
X_1588_ _0728_ _0732_ VGND VGND VPWR VPWR _0733_ sky130_fd_sc_hd__nor2_8
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2209_ _1088_ _1110_ _1236_ _1347_ _1348_ VGND VGND VPWR VPWR _1349_ sky130_fd_sc_hd__o221a_1
XFILLER_0_95_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2560_ _0206_ _0218_ _1197_ VGND VGND VPWR VPWR _0219_ sky130_fd_sc_hd__o21ai_1
X_2491_ _0136_ _0150_ VGND VGND VPWR VPWR _0151_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_50_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3112_ clknet_2_3__leaf_wb_clk_i _0007_ _0047_ VGND VGND VPWR VPWR weights_inst.data_out\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_77 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3043_ net14 net15 net16 VGND VGND VPWR VPWR _0690_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_77_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2827_ _1345_ _0813_ _1466_ _0483_ _1287_ VGND VGND VPWR VPWR _0485_ sky130_fd_sc_hd__o311a_1
XFILLER_0_60_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2758_ _1198_ _0408_ _0409_ _0411_ _0907_ VGND VGND VPWR VPWR _0412_ sky130_fd_sc_hd__a311o_1
XFILLER_0_60_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1709_ _0853_ VGND VGND VPWR VPWR _0854_ sky130_fd_sc_hd__clkbuf_8
X_2689_ _1232_ _1041_ _1025_ VGND VGND VPWR VPWR _0344_ sky130_fd_sc_hd__and3_1
XTAP_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1991_ _0667_ _1116_ _1122_ _1133_ _0860_ VGND VGND VPWR VPWR _1134_ sky130_fd_sc_hd__o311a_1
XFILLER_0_51_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2612_ _0263_ _0265_ _0268_ _1250_ _1164_ VGND VGND VPWR VPWR _0269_ sky130_fd_sc_hd__o221a_1
XFILLER_0_42_159 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2543_ _0962_ _1530_ _1140_ VGND VGND VPWR VPWR _0202_ sky130_fd_sc_hd__o21a_1
XFILLER_0_100_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2474_ _0861_ _1065_ _0093_ _0849_ VGND VGND VPWR VPWR _0135_ sky130_fd_sc_hd__a31o_1
XFILLER_0_76_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3026_ _0678_ VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__buf_1
XFILLER_0_93_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2190_ _1041_ _0976_ VGND VGND VPWR VPWR _1330_ sky130_fd_sc_hd__nor2_2
XFILLER_0_99_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1974_ _0745_ VGND VGND VPWR VPWR _1117_ sky130_fd_sc_hd__buf_4
XFILLER_0_70_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_498 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2526_ _1250_ _0179_ _0184_ _1273_ VGND VGND VPWR VPWR _0185_ sky130_fd_sc_hd__o211a_1
XFILLER_0_11_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2457_ _0936_ _0798_ _1112_ _0117_ _0934_ VGND VGND VPWR VPWR _0118_ sky130_fd_sc_hd__o311a_1
Xhold17 _1076_ VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__dlygate4sd3_1
Xhold28 net19 VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2388_ _0806_ _1020_ _1524_ _1060_ VGND VGND VPWR VPWR _1525_ sky130_fd_sc_hd__a211o_1
XFILLER_0_78_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3009_ weights_inst.data_out\[11\] _0666_ VGND VGND VPWR VPWR _0669_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1690_ _0834_ VGND VGND VPWR VPWR _0835_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_40_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2311_ _1052_ _1167_ VGND VGND VPWR VPWR _1449_ sky130_fd_sc_hd__nor2_2
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2242_ _1365_ _1378_ _1381_ _1322_ VGND VGND VPWR VPWR _1382_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_57_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2173_ _0735_ _0785_ VGND VGND VPWR VPWR _1314_ sky130_fd_sc_hd__nor2_4
XFILLER_0_73_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1957_ _0754_ _1099_ VGND VGND VPWR VPWR _1100_ sky130_fd_sc_hd__nor2_1
XFILLER_0_98_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1888_ _0763_ _1031_ VGND VGND VPWR VPWR _1032_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput29 net29 VGND VGND VPWR VPWR wbs_dat_o[18] sky130_fd_sc_hd__buf_12
X_2509_ _1198_ _0166_ _0168_ VGND VGND VPWR VPWR _0169_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_39_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_80 _1056_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2860_ _1396_ _0500_ _0507_ _0519_ VGND VGND VPWR VPWR _0520_ sky130_fd_sc_hd__o31a_1
XFILLER_0_84_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1811_ _0655_ _0850_ _0857_ _0859_ _0955_ VGND VGND VPWR VPWR _0004_ sky130_fd_sc_hd__o311a_1
XFILLER_0_65_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2791_ _0825_ _1015_ _0946_ _1236_ _0749_ VGND VGND VPWR VPWR _0446_ sky130_fd_sc_hd__a311o_1
XFILLER_0_53_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1742_ _0731_ _0886_ VGND VGND VPWR VPWR _0887_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_53_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1673_ _0717_ _0710_ VGND VGND VPWR VPWR _0818_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_25_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2225_ _1039_ VGND VGND VPWR VPWR _1365_ sky130_fd_sc_hd__buf_4
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2156_ _1273_ _1280_ _1286_ _1296_ _1161_ VGND VGND VPWR VPWR _1297_ sky130_fd_sc_hd__o311a_1
X_2087_ _1221_ VGND VGND VPWR VPWR _1229_ sky130_fd_sc_hd__buf_4
XFILLER_0_8_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2989_ net18 _0420_ _0657_ VGND VGND VPWR VPWR _0658_ sky130_fd_sc_hd__nor3_1
XFILLER_0_16_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2010_ _1140_ net52 _1150_ _1151_ _1152_ VGND VGND VPWR VPWR _1153_ sky130_fd_sc_hd__o32a_1
XFILLER_0_89_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2912_ _0575_ VGND VGND VPWR VPWR _0017_ sky130_fd_sc_hd__buf_1
XFILLER_0_57_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2843_ _0801_ _0977_ _1137_ _1043_ VGND VGND VPWR VPWR _0501_ sky130_fd_sc_hd__o22a_1
XFILLER_0_45_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2774_ _0900_ _0163_ _0427_ _0782_ VGND VGND VPWR VPWR _0428_ sky130_fd_sc_hd__o211a_1
X_1725_ _0718_ _0742_ _0741_ VGND VGND VPWR VPWR _0870_ sky130_fd_sc_hd__a21o_1
XFILLER_0_53_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1656_ _0800_ VGND VGND VPWR VPWR _0801_ sky130_fd_sc_hd__clkbuf_8
X_1587_ _0729_ _0731_ VGND VGND VPWR VPWR _0732_ sky130_fd_sc_hd__nand2_4
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2208_ _1056_ VGND VGND VPWR VPWR _1348_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_95_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2139_ _1274_ _1276_ _1277_ _1278_ _1279_ VGND VGND VPWR VPWR _1280_ sky130_fd_sc_hd__o311a_1
XFILLER_0_95_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2490_ _1243_ _0143_ _0149_ VGND VGND VPWR VPWR _0150_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_49_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3111_ clknet_2_2__leaf_wb_clk_i _0006_ _0046_ VGND VGND VPWR VPWR weights_inst.data_out\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_89 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3042_ net13 net14 net15 VGND VGND VPWR VPWR _0689_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_77_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2826_ _0873_ _1292_ _0266_ VGND VGND VPWR VPWR _0483_ sky130_fd_sc_hd__or3_1
XFILLER_0_45_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2757_ _1235_ _0966_ _1103_ _0410_ _0950_ VGND VGND VPWR VPWR _0411_ sky130_fd_sc_hd__o311a_1
XFILLER_0_76_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2688_ _0783_ _0337_ _0338_ _0342_ VGND VGND VPWR VPWR _0343_ sky130_fd_sc_hd__o31a_1
X_1708_ _0731_ _0759_ VGND VGND VPWR VPWR _0853_ sky130_fd_sc_hd__nand2_1
X_1639_ _0726_ VGND VGND VPWR VPWR _0784_ sky130_fd_sc_hd__buf_8
XTAP_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1990_ _1115_ _1126_ _1128_ _1132_ _0842_ VGND VGND VPWR VPWR _1133_ sky130_fd_sc_hd__a311o_1
XFILLER_0_67_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2611_ _1165_ _1206_ _1466_ _0267_ VGND VGND VPWR VPWR _0268_ sky130_fd_sc_hd__o31a_1
XFILLER_0_42_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2542_ _1219_ _1004_ _0890_ _0751_ VGND VGND VPWR VPWR _0201_ sky130_fd_sc_hd__a211o_2
XFILLER_0_2_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2473_ _0127_ _0133_ _1365_ VGND VGND VPWR VPWR _0134_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_76_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3025_ weights_inst.data_out\[19\] _0666_ VGND VGND VPWR VPWR _0678_ sky130_fd_sc_hd__and2_1
XFILLER_0_92_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2809_ _1403_ _1119_ _0273_ _0464_ _1308_ VGND VGND VPWR VPWR _0465_ sky130_fd_sc_hd__o311a_1
XFILLER_0_14_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1973_ _1109_ _1111_ _1112_ _1114_ _1115_ VGND VGND VPWR VPWR _1116_ sky130_fd_sc_hd__o311a_1
XFILLER_0_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2525_ _1047_ _0182_ _0183_ VGND VGND VPWR VPWR _0184_ sky130_fd_sc_hd__or3_1
X_2456_ _1136_ _0738_ _0929_ _1206_ _0956_ VGND VGND VPWR VPWR _0117_ sky130_fd_sc_hd__a221o_1
Xhold18 wbs_adr_i[6] VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__dlygate4sd3_1
X_2387_ _1015_ _0823_ _0738_ VGND VGND VPWR VPWR _1524_ sky130_fd_sc_hd__and3_2
XFILLER_0_78_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3008_ _0668_ VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__buf_1
XFILLER_0_78_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2310_ _1117_ _1097_ VGND VGND VPWR VPWR _1448_ sky130_fd_sc_hd__nor2_2
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2241_ _0892_ _1379_ _1380_ _1161_ VGND VGND VPWR VPWR _1381_ sky130_fd_sc_hd__a211o_1
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2172_ _0755_ _1232_ _1199_ _0805_ VGND VGND VPWR VPWR _1313_ sky130_fd_sc_hd__or4_1
XFILLER_0_28_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1956_ _0757_ _0767_ VGND VGND VPWR VPWR _1099_ sky130_fd_sc_hd__nor2_4
XFILLER_0_83_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1887_ _0795_ _0710_ VGND VGND VPWR VPWR _1031_ sky130_fd_sc_hd__nor2_4
XFILLER_0_101_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput19 net19 VGND VGND VPWR VPWR wbs_ack_o sky130_fd_sc_hd__buf_12
XFILLER_0_101_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2508_ _0931_ _1008_ _0167_ _0875_ _0914_ VGND VGND VPWR VPWR _0168_ sky130_fd_sc_hd__o221a_1
X_2439_ _0836_ _1045_ _1497_ VGND VGND VPWR VPWR _0100_ sky130_fd_sc_hd__or3b_1
XFILLER_0_94_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_70 _0764_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_81 _1063_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1810_ _0861_ _0909_ _0954_ VGND VGND VPWR VPWR _0955_ sky130_fd_sc_hd__or3_1
XFILLER_0_5_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2790_ _0910_ _1043_ _0444_ VGND VGND VPWR VPWR _0445_ sky130_fd_sc_hd__or3_1
XFILLER_0_13_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1741_ _0885_ VGND VGND VPWR VPWR _0886_ sky130_fd_sc_hd__buf_6
XFILLER_0_25_244 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1672_ _0765_ _0766_ VGND VGND VPWR VPWR _0817_ sky130_fd_sc_hd__nand2_8
XFILLER_0_53_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2224_ _0861_ _1333_ _1341_ _1353_ _1363_ VGND VGND VPWR VPWR _1364_ sky130_fd_sc_hd__o32a_1
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2155_ _1287_ _1290_ _1293_ _1295_ _0667_ VGND VGND VPWR VPWR _1296_ sky130_fd_sc_hd__a221o_1
XFILLER_0_76_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2086_ _1223_ _1227_ _0839_ VGND VGND VPWR VPWR _1228_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2988_ _0651_ _0656_ VGND VGND VPWR VPWR _0657_ sky130_fd_sc_hd__or2_1
XFILLER_0_44_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1939_ _1080_ _1081_ VGND VGND VPWR VPWR _1082_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2911_ net66 _0560_ _0574_ VGND VGND VPWR VPWR _0575_ sky130_fd_sc_hd__and3_1
XFILLER_0_73_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2842_ _0706_ _0496_ _0497_ _0499_ _1243_ VGND VGND VPWR VPWR _0500_ sky130_fd_sc_hd__a311oi_1
XFILLER_0_26_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2773_ _0964_ _1064_ _1475_ VGND VGND VPWR VPWR _0427_ sky130_fd_sc_hd__or3b_1
XFILLER_0_60_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1724_ _0852_ _0768_ VGND VGND VPWR VPWR _0869_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1655_ _0799_ VGND VGND VPWR VPWR _0800_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1586_ _0730_ VGND VGND VPWR VPWR _0731_ sky130_fd_sc_hd__buf_8
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2207_ _0786_ VGND VGND VPWR VPWR _1347_ sky130_fd_sc_hd__buf_4
XFILLER_0_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2138_ _0828_ _1084_ _1184_ _1264_ VGND VGND VPWR VPWR _1279_ sky130_fd_sc_hd__a211o_1
XFILLER_0_95_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2069_ _0835_ VGND VGND VPWR VPWR _1211_ sky130_fd_sc_hd__buf_4
XFILLER_0_76_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_49 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_158 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3110_ clknet_2_2__leaf_wb_clk_i _0005_ _0045_ VGND VGND VPWR VPWR weights_inst.data_out\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3041_ net13 VGND VGND VPWR VPWR _0688_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2825_ _1348_ _1044_ _1487_ _0481_ _0935_ VGND VGND VPWR VPWR _0482_ sky130_fd_sc_hd__o311a_1
XFILLER_0_14_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2756_ _0975_ _0976_ _1106_ _0802_ _0724_ VGND VGND VPWR VPWR _0410_ sky130_fd_sc_hd__a221o_1
XFILLER_0_14_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2687_ _0339_ _0341_ _0783_ VGND VGND VPWR VPWR _0342_ sky130_fd_sc_hd__o21ai_1
X_1707_ _0731_ _0737_ VGND VGND VPWR VPWR _0852_ sky130_fd_sc_hd__nand2_8
XFILLER_0_69_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1638_ _0782_ VGND VGND VPWR VPWR _0783_ sky130_fd_sc_hd__buf_4
X_1569_ net6 net4 VGND VGND VPWR VPWR _0714_ sky130_fd_sc_hd__nand2_2
XTAP_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2610_ _1030_ _0266_ _1165_ VGND VGND VPWR VPWR _0267_ sky130_fd_sc_hd__o21ai_1
X_2541_ _0762_ _1107_ VGND VGND VPWR VPWR _0200_ sky130_fd_sc_hd__or2b_1
X_2472_ _0706_ _0129_ _0132_ _0673_ VGND VGND VPWR VPWR _0133_ sky130_fd_sc_hd__a211o_1
XFILLER_0_11_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3024_ _0677_ VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__buf_1
XFILLER_0_92_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_158 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2808_ _1491_ _1016_ _0353_ VGND VGND VPWR VPWR _0464_ sky130_fd_sc_hd__or3_1
X_2739_ _0452_ _0813_ _0720_ VGND VGND VPWR VPWR _0393_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_41_194 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1972_ _0838_ VGND VGND VPWR VPWR _1115_ sky130_fd_sc_hd__buf_4
XFILLER_0_28_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2524_ _1056_ _0893_ _1456_ VGND VGND VPWR VPWR _0183_ sky130_fd_sc_hd__nor3_1
XFILLER_0_11_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2455_ _0086_ _0115_ _0764_ VGND VGND VPWR VPWR _0116_ sky130_fd_sc_hd__a21o_1
Xhold19 _0846_ VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__dlygate4sd3_1
X_2386_ _0852_ _0970_ _1025_ VGND VGND VPWR VPWR _1523_ sky130_fd_sc_hd__and3_1
XFILLER_0_78_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3007_ weights_inst.data_out\[10\] _0666_ VGND VGND VPWR VPWR _0668_ sky130_fd_sc_hd__and2_1
XFILLER_0_93_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2240_ _0758_ _0831_ _0947_ VGND VGND VPWR VPWR _1380_ sky130_fd_sc_hd__and3_2
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2171_ _1311_ _1064_ _1190_ _0945_ _0977_ VGND VGND VPWR VPWR _1312_ sky130_fd_sc_hd__a221o_1
XFILLER_0_73_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1955_ _0769_ _1097_ VGND VGND VPWR VPWR _1098_ sky130_fd_sc_hd__nand2_2
XFILLER_0_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1886_ _0745_ _0760_ VGND VGND VPWR VPWR _1030_ sky130_fd_sc_hd__nor2_4
XFILLER_0_43_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2507_ _1113_ _0744_ _0948_ VGND VGND VPWR VPWR _0167_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_51_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2438_ _1335_ _1248_ _0098_ VGND VGND VPWR VPWR _0099_ sky130_fd_sc_hd__mux2_1
X_2369_ _0892_ _0973_ VGND VGND VPWR VPWR _1506_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_71 _0782_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_82 _1064_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_60 _1407_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_cap51 _1422_ VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__buf_2
XFILLER_0_97_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1740_ _0717_ net3 VGND VGND VPWR VPWR _0885_ sky130_fd_sc_hd__and2_1
XFILLER_0_25_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1671_ _0815_ VGND VGND VPWR VPWR _0816_ sky130_fd_sc_hd__buf_4
XFILLER_0_13_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2223_ _1273_ _1357_ _1362_ _0645_ VGND VGND VPWR VPWR _1363_ sky130_fd_sc_hd__a31o_1
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2154_ _0971_ _1079_ _1294_ _0751_ VGND VGND VPWR VPWR _1295_ sky130_fd_sc_hd__a211o_1
X_2085_ _1044_ _1225_ _1226_ VGND VGND VPWR VPWR _1227_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_76_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2987_ net6 net4 net7 net5 VGND VGND VPWR VPWR _0656_ sky130_fd_sc_hd__or4_1
X_1938_ _0916_ _1045_ _0912_ _0724_ VGND VGND VPWR VPWR _1081_ sky130_fd_sc_hd__a211o_1
XFILLER_0_71_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1869_ _0823_ VGND VGND VPWR VPWR _1013_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_44_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2910_ _0645_ _0572_ _0573_ _1497_ _0848_ VGND VGND VPWR VPWR _0574_ sky130_fd_sc_hd__a221o_1
XFILLER_0_57_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2841_ _1252_ _0316_ _0498_ _0935_ VGND VGND VPWR VPWR _0499_ sky130_fd_sc_hd__o211a_1
XFILLER_0_57_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2772_ _0952_ _0416_ _0419_ _0425_ _0860_ VGND VGND VPWR VPWR _0426_ sky130_fd_sc_hd__o311a_1
XFILLER_0_13_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1723_ _0708_ _0765_ VGND VGND VPWR VPWR _0868_ sky130_fd_sc_hd__nor2_8
X_1654_ _0723_ VGND VGND VPWR VPWR _0799_ sky130_fd_sc_hd__buf_4
X_1585_ net6 net4 VGND VGND VPWR VPWR _0730_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_21_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2206_ _1343_ _0868_ _1344_ _1345_ VGND VGND VPWR VPWR _1346_ sky130_fd_sc_hd__o211a_1
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2137_ _0950_ VGND VGND VPWR VPWR _1278_ sky130_fd_sc_hd__buf_4
X_2068_ _0881_ _0800_ _0805_ _1077_ VGND VGND VPWR VPWR _1210_ sky130_fd_sc_hd__or4_1
XFILLER_0_76_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3040_ _0687_ VGND VGND VPWR VPWR _0002_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2824_ _1000_ _1229_ _0819_ _1199_ _1109_ VGND VGND VPWR VPWR _0481_ sky130_fd_sc_hd__a221o_1
XFILLER_0_14_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2755_ _0865_ _1184_ VGND VGND VPWR VPWR _0409_ sky130_fd_sc_hd__or2_1
X_2686_ _0852_ _1311_ _0340_ _1300_ _0923_ VGND VGND VPWR VPWR _0341_ sky130_fd_sc_hd__o221a_1
X_1706_ _0729_ _0735_ VGND VGND VPWR VPWR _0851_ sky130_fd_sc_hd__nand2_4
XFILLER_0_1_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1637_ _0777_ VGND VGND VPWR VPWR _0782_ sky130_fd_sc_hd__clkbuf_8
XTAP_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1568_ _0712_ VGND VGND VPWR VPWR _0713_ sky130_fd_sc_hd__buf_4
XTAP_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2540_ _1348_ _1129_ _0124_ _0198_ _1285_ VGND VGND VPWR VPWR _0199_ sky130_fd_sc_hd__o311a_1
X_2471_ _1348_ _0774_ _1059_ _0131_ _0779_ VGND VGND VPWR VPWR _0132_ sky130_fd_sc_hd__o311a_1
X_3023_ weights_inst.data_out\[18\] _0666_ VGND VGND VPWR VPWR _0677_ sky130_fd_sc_hd__and2_1
XFILLER_0_18_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2807_ _0460_ _0344_ _0461_ _1285_ VGND VGND VPWR VPWR _0463_ sky130_fd_sc_hd__o211a_1
X_2738_ _1281_ _0807_ _0389_ _0391_ _1285_ VGND VGND VPWR VPWR _0392_ sky130_fd_sc_hd__o311a_1
XFILLER_0_41_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2669_ _1000_ _0917_ _0819_ _1311_ _1180_ VGND VGND VPWR VPWR _0325_ sky130_fd_sc_hd__a221o_1
XFILLER_0_1_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1971_ _1113_ _1072_ _0929_ _0925_ _0750_ VGND VGND VPWR VPWR _1114_ sky130_fd_sc_hd__a221o_1
XFILLER_0_83_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2523_ _0743_ _1188_ _0181_ _0810_ VGND VGND VPWR VPWR _0182_ sky130_fd_sc_hd__o211a_1
XFILLER_0_23_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2454_ _1019_ _0855_ _1060_ VGND VGND VPWR VPWR _0115_ sky130_fd_sc_hd__a21o_1
X_2385_ _0803_ _0816_ _1030_ _0735_ _1040_ VGND VGND VPWR VPWR _1522_ sky130_fd_sc_hd__a221o_1
Xinput1 wb_rst_i VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_2
X_3006_ net55 VGND VGND VPWR VPWR _0666_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_93_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2170_ _0970_ VGND VGND VPWR VPWR _1311_ sky130_fd_sc_hd__buf_4
XFILLER_0_73_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1954_ _0891_ _0973_ _0886_ VGND VGND VPWR VPWR _1097_ sky130_fd_sc_hd__a21o_4
XFILLER_0_28_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1885_ _1026_ _1027_ _1028_ VGND VGND VPWR VPWR _1029_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_98_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2506_ _0725_ _0163_ _0164_ _0165_ VGND VGND VPWR VPWR _0166_ sky130_fd_sc_hd__o31a_1
X_2437_ _0871_ _1360_ VGND VGND VPWR VPWR _0098_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2368_ _1311_ net52 _1026_ _1040_ VGND VGND VPWR VPWR _1505_ sky130_fd_sc_hd__a211o_1
XFILLER_0_98_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2299_ _0810_ _1103_ _1302_ _1436_ _0694_ VGND VGND VPWR VPWR _1437_ sky130_fd_sc_hd__o311a_1
XFILLER_0_78_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_50 _1160_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_72 _0782_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_83 _1190_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_61 _1407_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1670_ _0814_ VGND VGND VPWR VPWR _0815_ sky130_fd_sc_hd__buf_4
XFILLER_0_40_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2222_ _1274_ _1358_ _1359_ _1361_ _1178_ VGND VGND VPWR VPWR _1362_ sky130_fd_sc_hd__a311o_1
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2153_ _1015_ _0887_ VGND VGND VPWR VPWR _1294_ sky130_fd_sc_hd__and2_4
X_2084_ _1184_ _0724_ _1055_ VGND VGND VPWR VPWR _1226_ sky130_fd_sc_hd__or3b_1
XFILLER_0_75_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_94 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2986_ _0653_ VGND VGND VPWR VPWR _0654_ sky130_fd_sc_hd__buf_2
XFILLER_0_29_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1937_ _0983_ _1077_ _1079_ _0971_ _0910_ VGND VGND VPWR VPWR _1080_ sky130_fd_sc_hd__a221o_1
XFILLER_0_71_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1868_ _0852_ _1003_ VGND VGND VPWR VPWR _1012_ sky130_fd_sc_hd__nand2_2
XFILLER_0_101_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1799_ _0834_ VGND VGND VPWR VPWR _0944_ sky130_fd_sc_hd__buf_4
XFILLER_0_79_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2840_ _1063_ _1249_ _0467_ VGND VGND VPWR VPWR _0498_ sky130_fd_sc_hd__or3_1
XFILLER_0_57_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_382 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2771_ _1115_ _0421_ _0422_ _0424_ _0993_ VGND VGND VPWR VPWR _0425_ sky130_fd_sc_hd__a311o_1
XFILLER_0_13_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1722_ _0866_ VGND VGND VPWR VPWR _0867_ sky130_fd_sc_hd__buf_4
XFILLER_0_79_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1653_ _0794_ _0728_ _0797_ VGND VGND VPWR VPWR _0798_ sky130_fd_sc_hd__and3_4
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1584_ net3 VGND VGND VPWR VPWR _0729_ sky130_fd_sc_hd__inv_6
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2205_ _0936_ VGND VGND VPWR VPWR _1345_ sky130_fd_sc_hd__clkbuf_4
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2136_ _0716_ _0866_ _0959_ VGND VGND VPWR VPWR _1277_ sky130_fd_sc_hd__and3_4
X_2067_ _1198_ _1201_ _1203_ _1208_ VGND VGND VPWR VPWR _1209_ sky130_fd_sc_hd__a31o_1
XFILLER_0_44_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2969_ _0633_ _0636_ _1243_ VGND VGND VPWR VPWR _0637_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_71_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_308 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2823_ _0459_ _0466_ _0479_ VGND VGND VPWR VPWR _0480_ sky130_fd_sc_hd__a21oi_1
X_2754_ _1219_ _1004_ _1084_ _1056_ VGND VGND VPWR VPWR _0408_ sky130_fd_sc_hd__a211o_1
XFILLER_0_26_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1705_ _0673_ _0781_ _0844_ _0849_ VGND VGND VPWR VPWR _0850_ sky130_fd_sc_hd__o211a_1
XFILLER_0_41_311 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2685_ _0756_ _0760_ VGND VGND VPWR VPWR _0340_ sky130_fd_sc_hd__nor2_4
X_1636_ _0706_ _0753_ _0780_ VGND VGND VPWR VPWR _0781_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1567_ _0708_ _0711_ VGND VGND VPWR VPWR _0712_ sky130_fd_sc_hd__nand2_4
XTAP_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2119_ _1019_ _1043_ _1259_ VGND VGND VPWR VPWR _1260_ sky130_fd_sc_hd__a21o_1
X_3099_ clknet_2_1__leaf_wb_clk_i net86 _0034_ VGND VGND VPWR VPWR fsm_inst.current_state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2470_ _1211_ _1418_ _0130_ VGND VGND VPWR VPWR _0131_ sky130_fd_sc_hd__or3_1
XFILLER_0_50_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3022_ _0676_ VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__buf_1
XFILLER_0_19_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2806_ _0873_ _1491_ _1463_ VGND VGND VPWR VPWR _0461_ sky130_fd_sc_hd__or3_1
X_2737_ _0390_ _0983_ _1261_ VGND VGND VPWR VPWR _0391_ sky130_fd_sc_hd__a21o_1
XFILLER_0_74_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2668_ _1273_ _0315_ _0318_ _0323_ _1161_ VGND VGND VPWR VPWR _0324_ sky130_fd_sc_hd__o311a_1
X_1619_ _0763_ _0719_ _0712_ VGND VGND VPWR VPWR _0764_ sky130_fd_sc_hd__and3_4
X_2599_ _0878_ _0989_ VGND VGND VPWR VPWR _0256_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_360 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1970_ _0735_ _0999_ VGND VGND VPWR VPWR _1113_ sky130_fd_sc_hd__nand2_2
XFILLER_0_95_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_299 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2522_ _0970_ _0180_ VGND VGND VPWR VPWR _0181_ sky130_fd_sc_hd__nand2_2
XFILLER_0_87_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2453_ _1023_ _1253_ _0113_ _1135_ _1198_ VGND VGND VPWR VPWR _0114_ sky130_fd_sc_hd__o221a_1
X_2384_ _1335_ _1519_ _1520_ VGND VGND VPWR VPWR _1521_ sky130_fd_sc_hd__nand3_1
Xinput2 net79 VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_2
X_3005_ _0665_ VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__buf_1
XFILLER_0_36_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_494 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1953_ _0724_ _1095_ VGND VGND VPWR VPWR _1096_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1884_ _0834_ VGND VGND VPWR VPWR _1028_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_28_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_450 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2505_ _0984_ _0999_ _0814_ _1491_ VGND VGND VPWR VPWR _0165_ sky130_fd_sc_hd__or4_1
X_2436_ _1158_ _0067_ _0068_ _0859_ _0097_ VGND VGND VPWR VPWR _0027_ sky130_fd_sc_hd__o311a_1
XFILLER_0_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2367_ _1311_ _0867_ _0892_ _1379_ _1180_ VGND VGND VPWR VPWR _1504_ sky130_fd_sc_hd__a221o_1
X_2298_ _0806_ _1020_ _1097_ _1117_ _0835_ VGND VGND VPWR VPWR _1436_ sky130_fd_sc_hd__a221o_1
XFILLER_0_78_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_40 _1038_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_73 _0798_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_62 _1407_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_84 _1190_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_51 _1173_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap53 _0658_ VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__buf_1
XFILLER_0_85_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2221_ _0919_ _1360_ _1261_ VGND VGND VPWR VPWR _1361_ sky130_fd_sc_hd__a21oi_1
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2152_ _1291_ _1292_ _0703_ VGND VGND VPWR VPWR _1293_ sky130_fd_sc_hd__a21oi_1
X_2083_ _0834_ _1224_ VGND VGND VPWR VPWR _1225_ sky130_fd_sc_hd__or2_2
XFILLER_0_88_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2985_ net18 _0420_ _0651_ _0652_ VGND VGND VPWR VPWR _0653_ sky130_fd_sc_hd__nor4_1
XFILLER_0_29_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1936_ _0939_ _1078_ VGND VGND VPWR VPWR _1079_ sky130_fd_sc_hd__nor2_4
X_1867_ _0785_ VGND VGND VPWR VPWR _1011_ sky130_fd_sc_hd__buf_4
XFILLER_0_44_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1798_ _0936_ _0938_ _0940_ net52 _0942_ VGND VGND VPWR VPWR _0943_ sky130_fd_sc_hd__o32a_1
XFILLER_0_12_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2419_ _1090_ _0080_ _0984_ VGND VGND VPWR VPWR _0081_ sky130_fd_sc_hd__and3b_1
XFILLER_0_94_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2770_ _0944_ _0940_ _1079_ _0423_ _0777_ VGND VGND VPWR VPWR _0424_ sky130_fd_sc_hd__o311a_2
XFILLER_0_38_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1721_ _0729_ _0711_ VGND VGND VPWR VPWR _0866_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_26_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1652_ _0796_ VGND VGND VPWR VPWR _0797_ sky130_fd_sc_hd__buf_4
XFILLER_0_0_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1583_ _0727_ VGND VGND VPWR VPWR _0728_ sky130_fd_sc_hd__buf_8
XFILLER_0_95_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2204_ _0867_ _1030_ VGND VGND VPWR VPWR _1344_ sky130_fd_sc_hd__nand2_1
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2135_ _0760_ _1275_ VGND VGND VPWR VPWR _1276_ sky130_fd_sc_hd__nor2_2
XFILLER_0_76_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2066_ _0875_ _1206_ _1094_ _1207_ _0950_ VGND VGND VPWR VPWR _1208_ sky130_fd_sc_hd__o311a_1
XFILLER_0_48_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2968_ _0595_ _0635_ _0783_ VGND VGND VPWR VPWR _0636_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_71_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1919_ _0754_ VGND VGND VPWR VPWR _1063_ sky130_fd_sc_hd__buf_8
XFILLER_0_60_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2899_ _0964_ _0941_ _1230_ _0561_ _0913_ VGND VGND VPWR VPWR _0562_ sky130_fd_sc_hd__o32a_1
XFILLER_0_44_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2822_ _0673_ _0469_ _0471_ _0478_ _1396_ VGND VGND VPWR VPWR _0479_ sky130_fd_sc_hd__o311a_1
XFILLER_0_38_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2753_ _1278_ _0403_ _0404_ _0406_ _1193_ VGND VGND VPWR VPWR _0407_ sky130_fd_sc_hd__a311o_1
X_1704_ _0848_ VGND VGND VPWR VPWR _0849_ sky130_fd_sc_hd__buf_8
XFILLER_0_41_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2684_ _1067_ _1519_ _1291_ VGND VGND VPWR VPWR _0339_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1635_ _0762_ _0764_ _0775_ _0752_ _0779_ VGND VGND VPWR VPWR _0780_ sky130_fd_sc_hd__o221a_1
XFILLER_0_22_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1566_ _0710_ VGND VGND VPWR VPWR _0711_ sky130_fd_sc_hd__buf_12
XTAP_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3098_ clknet_2_1__leaf_wb_clk_i net63 _0033_ VGND VGND VPWR VPWR fsm_inst.current_state\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_2118_ _0786_ _0788_ _1063_ VGND VGND VPWR VPWR _1259_ sky130_fd_sc_hd__o21ai_4
X_2049_ _0980_ _1190_ VGND VGND VPWR VPWR _1191_ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3021_ weights_inst.data_out\[17\] _0666_ VGND VGND VPWR VPWR _0676_ sky130_fd_sc_hd__and2_1
XFILLER_0_18_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2805_ _1274_ _0919_ VGND VGND VPWR VPWR _0460_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2736_ _0806_ _0867_ VGND VGND VPWR VPWR _0390_ sky130_fd_sc_hd__nand2_1
X_2667_ _1287_ _0319_ _0320_ _0322_ _0667_ VGND VGND VPWR VPWR _0323_ sky130_fd_sc_hd__a311o_1
XFILLER_0_67_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1618_ _0715_ VGND VGND VPWR VPWR _0763_ sky130_fd_sc_hd__clkbuf_4
X_2598_ _1158_ _0232_ _0255_ _1242_ VGND VGND VPWR VPWR _0008_ sky130_fd_sc_hd__o211a_1
X_1549_ _0516_ _0580_ VGND VGND VPWR VPWR _0591_ sky130_fd_sc_hd__and2_1
XTAP_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2521_ _1089_ _0867_ VGND VGND VPWR VPWR _0180_ sky130_fd_sc_hd__nand2_2
XFILLER_0_11_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2452_ _1235_ _1294_ VGND VGND VPWR VPWR _0113_ sky130_fd_sc_hd__or2_1
X_2383_ _1043_ _0916_ VGND VGND VPWR VPWR _1520_ sky130_fd_sc_hd__nand2_1
X_3004_ weights_inst.data_out\[9\] _0654_ VGND VGND VPWR VPWR _0665_ sky130_fd_sc_hd__and2_1
Xinput3 net73 VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__buf_4
XFILLER_0_93_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2719_ _0634_ _0371_ _0373_ VGND VGND VPWR VPWR _0374_ sky130_fd_sc_hd__or3_1
XFILLER_0_30_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1952_ _0802_ _1072_ VGND VGND VPWR VPWR _1095_ sky130_fd_sc_hd__nand2_1
XFILLER_0_83_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1883_ _0763_ _0796_ _0946_ VGND VGND VPWR VPWR _1027_ sky130_fd_sc_hd__and3_2
XFILLER_0_56_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2504_ _1117_ _0976_ _1073_ VGND VGND VPWR VPWR _0164_ sky130_fd_sc_hd__and3_1
XFILLER_0_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2435_ _0863_ _0084_ _0096_ VGND VGND VPWR VPWR _0097_ sky130_fd_sc_hd__or3_1
XFILLER_0_47_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2366_ _1403_ _1500_ _1501_ _0935_ _1502_ VGND VGND VPWR VPWR _1503_ sky130_fd_sc_hd__o311a_1
X_2297_ _1140_ _1432_ _1433_ _1434_ _0694_ VGND VGND VPWR VPWR _1435_ sky130_fd_sc_hd__o311a_1
XFILLER_0_47_83 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_41 _1038_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_30 _0898_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_52 _1200_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_63 _1407_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_74 _0798_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_85 _1265_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmax_cap54 _0880_ VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__buf_4
XFILLER_0_69_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2220_ _1003_ _0770_ VGND VGND VPWR VPWR _1360_ sky130_fd_sc_hd__nand2_1
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2151_ _0881_ _0819_ _0820_ VGND VGND VPWR VPWR _1292_ sky130_fd_sc_hd__a21oi_2
X_2082_ _0828_ _0763_ _0866_ VGND VGND VPWR VPWR _1224_ sky130_fd_sc_hd__and3_1
XFILLER_0_88_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2984_ net6 net4 net7 net5 VGND VGND VPWR VPWR _0652_ sky130_fd_sc_hd__or4b_1
XFILLER_0_44_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1935_ net57 VGND VGND VPWR VPWR _1078_ sky130_fd_sc_hd__buf_6
XFILLER_0_83_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1866_ _1008_ _1009_ VGND VGND VPWR VPWR _1010_ sky130_fd_sc_hd__or2_1
X_1797_ _0754_ _0941_ VGND VGND VPWR VPWR _0942_ sky130_fd_sc_hd__or2_2
XFILLER_0_58_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2418_ _0831_ _0892_ _0973_ _0740_ VGND VGND VPWR VPWR _0080_ sky130_fd_sc_hd__a31o_2
XFILLER_0_58_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2349_ _1244_ _0733_ _0813_ _1485_ _1342_ VGND VGND VPWR VPWR _1486_ sky130_fd_sc_hd__o311a_1
XFILLER_0_94_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1720_ _0825_ _0769_ _0864_ VGND VGND VPWR VPWR _0865_ sky130_fd_sc_hd__a21o_1
XFILLER_0_41_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1651_ _0795_ _0731_ VGND VGND VPWR VPWR _0796_ sky130_fd_sc_hd__nand2_2
X_1582_ _0726_ VGND VGND VPWR VPWR _0727_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_0_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2203_ _0878_ VGND VGND VPWR VPWR _1343_ sky130_fd_sc_hd__clkbuf_4
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2134_ _0745_ _0712_ VGND VGND VPWR VPWR _1275_ sky130_fd_sc_hd__nand2_4
XFILLER_0_88_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2065_ _0803_ _0815_ _1137_ _0964_ VGND VGND VPWR VPWR _1207_ sky130_fd_sc_hd__a211o_1
XFILLER_0_76_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2967_ _0110_ _0186_ _1256_ VGND VGND VPWR VPWR _0635_ sky130_fd_sc_hd__a21o_1
XFILLER_0_8_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1918_ _1000_ _1043_ _1016_ _0890_ _0800_ VGND VGND VPWR VPWR _1062_ sky130_fd_sc_hd__a2111o_1
X_2898_ _0785_ _0380_ _0749_ VGND VGND VPWR VPWR _0561_ sky130_fd_sc_hd__a21o_1
XFILLER_0_44_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1849_ _0661_ VGND VGND VPWR VPWR _0993_ sky130_fd_sc_hd__buf_4
XFILLER_0_69_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2821_ _1342_ _0475_ _0477_ _0952_ VGND VGND VPWR VPWR _0478_ sky130_fd_sc_hd__a211o_1
XFILLER_0_26_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2752_ _0923_ _1392_ _1520_ _0405_ _1115_ VGND VGND VPWR VPWR _0406_ sky130_fd_sc_hd__a311oi_1
XFILLER_0_38_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1703_ _0845_ net78 net69 VGND VGND VPWR VPWR _0848_ sky130_fd_sc_hd__nand3_4
XFILLER_0_26_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2683_ _0771_ _1347_ _0760_ _1453_ _1274_ VGND VGND VPWR VPWR _0338_ sky130_fd_sc_hd__o311a_1
XFILLER_0_41_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1634_ _0778_ VGND VGND VPWR VPWR _0779_ sky130_fd_sc_hd__clkbuf_4
X_1565_ net6 net4 VGND VGND VPWR VPWR _0710_ sky130_fd_sc_hd__xor2_4
XTAP_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3097_ clknet_2_1__leaf_wb_clk_i net61 _0032_ VGND VGND VPWR VPWR fsm_inst.current_state\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_2117_ _1183_ _1253_ _1257_ _0706_ VGND VGND VPWR VPWR _1258_ sky130_fd_sc_hd__o211a_1
X_2048_ _0825_ _0877_ VGND VGND VPWR VPWR _1190_ sky130_fd_sc_hd__nor2_8
XFILLER_0_12_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_107 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3020_ _0675_ VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__buf_1
XFILLER_0_25_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_86 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2804_ _1164_ _0456_ _0458_ VGND VGND VPWR VPWR _0459_ sky130_fd_sc_hd__or3_1
XFILLER_0_73_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2735_ _1123_ _0877_ VGND VGND VPWR VPWR _0389_ sky130_fd_sc_hd__nor2_2
X_2666_ _1056_ _0903_ _1379_ _0321_ _0778_ VGND VGND VPWR VPWR _0322_ sky130_fd_sc_hd__o311a_1
X_1617_ _0755_ _0761_ VGND VGND VPWR VPWR _0762_ sky130_fd_sc_hd__nand2_1
X_2597_ _1365_ _0242_ _0254_ _1322_ VGND VGND VPWR VPWR _0255_ sky130_fd_sc_hd__a211o_1
X_1548_ _0548_ _0570_ VGND VGND VPWR VPWR _0580_ sky130_fd_sc_hd__xnor2_4
XTAP_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_419 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2520_ _1343_ _0819_ _0976_ _0811_ _0737_ VGND VGND VPWR VPWR _0179_ sky130_fd_sc_hd__a221o_1
XFILLER_0_11_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_474 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2451_ _1256_ _1282_ _0109_ _0111_ _1278_ VGND VGND VPWR VPWR _0112_ sky130_fd_sc_hd__o311a_1
X_2382_ _0807_ _0976_ VGND VGND VPWR VPWR _1519_ sky130_fd_sc_hd__nand2_1
Xinput4 net81 VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__buf_4
X_3003_ _0664_ VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__buf_1
XFILLER_0_59_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2718_ _1109_ _0902_ _0372_ _0963_ VGND VGND VPWR VPWR _0373_ sky130_fd_sc_hd__o211a_1
XFILLER_0_14_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2649_ _1147_ _0303_ _0304_ _0935_ VGND VGND VPWR VPWR _0305_ sky130_fd_sc_hd__o211a_1
XFILLER_0_100_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1951_ _0939_ _0713_ _0892_ VGND VGND VPWR VPWR _1094_ sky130_fd_sc_hd__and3_2
XFILLER_0_83_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1882_ _0740_ _0796_ _1025_ VGND VGND VPWR VPWR _1026_ sky130_fd_sc_hd__and3_2
X_2503_ _1041_ _1013_ _0738_ VGND VGND VPWR VPWR _0163_ sky130_fd_sc_hd__and3_1
XFILLER_0_11_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2434_ _0843_ _0087_ _0090_ _0095_ _0645_ VGND VGND VPWR VPWR _0096_ sky130_fd_sc_hd__o311a_1
X_2365_ _0936_ _0988_ _1200_ VGND VGND VPWR VPWR _1502_ sky130_fd_sc_hd__or3_1
X_2296_ _1305_ _0749_ _0961_ VGND VGND VPWR VPWR _1434_ sky130_fd_sc_hd__or3b_1
XFILLER_0_47_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_83 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_31 _0900_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_20 _0725_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_42 _1038_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_75 _0898_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_64 _1470_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_53 _1200_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_86 _1399_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_308 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2150_ _1063_ VGND VGND VPWR VPWR _1291_ sky130_fd_sc_hd__buf_4
X_2081_ _1019_ _1219_ _1220_ _1222_ _1211_ VGND VGND VPWR VPWR _1223_ sky130_fd_sc_hd__a32o_1
XFILLER_0_88_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_87 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2983_ net8 net9 net10 net85 VGND VGND VPWR VPWR _0651_ sky130_fd_sc_hd__or4_1
X_1934_ _0757_ _0901_ VGND VGND VPWR VPWR _1077_ sky130_fd_sc_hd__nor2_4
XFILLER_0_83_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1865_ _0877_ _0738_ _0817_ VGND VGND VPWR VPWR _1009_ sky130_fd_sc_hd__and3_1
XFILLER_0_44_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1796_ _0758_ _0866_ VGND VGND VPWR VPWR _0941_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2417_ _0820_ _0738_ _0937_ _1325_ VGND VGND VPWR VPWR _0079_ sky130_fd_sc_hd__a31o_1
XFILLER_0_42_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2348_ _1073_ _1379_ _1439_ _0923_ VGND VGND VPWR VPWR _1485_ sky130_fd_sc_hd__a211o_1
X_2279_ _0881_ _0918_ _0797_ VGND VGND VPWR VPWR _1418_ sky130_fd_sc_hd__and3_1
XFILLER_0_67_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1650_ net2 VGND VGND VPWR VPWR _0795_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1581_ net58 _0714_ VGND VGND VPWR VPWR _0726_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_1_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2202_ _1115_ VGND VGND VPWR VPWR _1342_ sky130_fd_sc_hd__buf_4
X_2133_ _0875_ VGND VGND VPWR VPWR _1274_ sky130_fd_sc_hd__buf_4
X_2064_ _1205_ VGND VGND VPWR VPWR _1206_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_44_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2966_ _1335_ _0721_ _0590_ _0632_ _0935_ VGND VGND VPWR VPWR _0633_ sky130_fd_sc_hd__o311a_1
X_1917_ _0946_ _1059_ _1060_ _0832_ VGND VGND VPWR VPWR _1061_ sky130_fd_sc_hd__a211o_1
X_2897_ _0545_ _0558_ _0849_ VGND VGND VPWR VPWR _0560_ sky130_fd_sc_hd__o21ai_4
X_1848_ _0750_ _0925_ _0988_ _0991_ _0838_ VGND VGND VPWR VPWR _0992_ sky130_fd_sc_hd__o311a_1
XFILLER_0_8_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1779_ _0746_ VGND VGND VPWR VPWR _0924_ sky130_fd_sc_hd__buf_4
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2820_ _0751_ _1418_ _1449_ _0476_ _0782_ VGND VGND VPWR VPWR _0477_ sky130_fd_sc_hd__o311a_1
XFILLER_0_26_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2751_ _0786_ _0929_ _1174_ _1063_ VGND VGND VPWR VPWR _0405_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_81_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1702_ _0613_ net10 net9 VGND VGND VPWR VPWR _0847_ sky130_fd_sc_hd__nand3b_1
X_2682_ _0900_ _1003_ VGND VGND VPWR VPWR _0337_ sky130_fd_sc_hd__and2b_1
XFILLER_0_26_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1633_ _0777_ VGND VGND VPWR VPWR _0778_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_30_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1564_ net3 VGND VGND VPWR VPWR _0708_ sky130_fd_sc_hd__buf_8
XTAP_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3096_ clknet_2_1__leaf_wb_clk_i _0000_ _0031_ VGND VGND VPWR VPWR fsm_inst.cnn_en
+ sky130_fd_sc_hd__dfrtp_1
X_2116_ _1124_ _0816_ _1255_ _1256_ VGND VGND VPWR VPWR _1257_ sky130_fd_sc_hd__a211o_1
XFILLER_0_89_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2047_ _1188_ net56 VGND VGND VPWR VPWR _1189_ sky130_fd_sc_hd__nor2_2
XFILLER_0_76_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2949_ _0723_ _0764_ _0888_ VGND VGND VPWR VPWR _0616_ sky130_fd_sc_hd__or3_1
XFILLER_0_17_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_244 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2803_ _1345_ _0855_ _1213_ _0457_ _1287_ VGND VGND VPWR VPWR _0458_ sky130_fd_sc_hd__o311a_1
XFILLER_0_41_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2734_ _0673_ _0379_ _0382_ _0387_ _0655_ VGND VGND VPWR VPWR _0388_ sky130_fd_sc_hd__o311a_1
XFILLER_0_41_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2665_ _0835_ _0733_ _0855_ VGND VGND VPWR VPWR _0321_ sky130_fd_sc_hd__or3_1
X_2596_ _0861_ _0253_ VGND VGND VPWR VPWR _0254_ sky130_fd_sc_hd__nor2_1
X_1616_ _0756_ _0758_ _0760_ VGND VGND VPWR VPWR _0761_ sky130_fd_sc_hd__or3_4
XFILLER_0_10_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1547_ net6 net8 _0441_ _0559_ VGND VGND VPWR VPWR _0570_ sky130_fd_sc_hd__a31o_2
XFILLER_0_66_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3079_ _0707_ VGND VGND VPWR VPWR _0046_ sky130_fd_sc_hd__inv_2
XFILLER_0_92_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_255 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_450 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_306 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2450_ _1275_ _0110_ _0751_ VGND VGND VPWR VPWR _0111_ sky130_fd_sc_hd__a21o_1
XFILLER_0_51_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2381_ _1515_ _1517_ _0706_ VGND VGND VPWR VPWR _1518_ sky130_fd_sc_hd__a21oi_1
Xinput5 net83 VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_2
X_3002_ weights_inst.data_out\[8\] _0654_ VGND VGND VPWR VPWR _0664_ sky130_fd_sc_hd__and2_1
XFILLER_0_59_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_388 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2717_ _0916_ _1152_ _0266_ _0750_ VGND VGND VPWR VPWR _0372_ sky130_fd_sc_hd__a211o_1
XFILLER_0_72_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2648_ _1235_ _1380_ _1511_ VGND VGND VPWR VPWR _0304_ sky130_fd_sc_hd__or3_1
X_2579_ _0760_ _0867_ VGND VGND VPWR VPWR _0237_ sky130_fd_sc_hd__nor2_1
XFILLER_0_100_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1950_ _0964_ _0760_ _1088_ _1059_ _1092_ VGND VGND VPWR VPWR _1093_ sky130_fd_sc_hd__o41a_1
XFILLER_0_56_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1881_ _0735_ _0760_ VGND VGND VPWR VPWR _1025_ sky130_fd_sc_hd__nand2_4
XFILLER_0_56_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_250 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2502_ _1178_ _0158_ _0159_ _0161_ VGND VGND VPWR VPWR _0162_ sky130_fd_sc_hd__a31o_1
XFILLER_0_11_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2433_ _0839_ _0092_ _0094_ _1098_ _0907_ VGND VGND VPWR VPWR _0095_ sky130_fd_sc_hd__a221o_1
X_2364_ _0770_ _0788_ VGND VGND VPWR VPWR _1501_ sky130_fd_sc_hd__nor2_1
X_2295_ _0772_ _0926_ _1391_ VGND VGND VPWR VPWR _1433_ sky130_fd_sc_hd__and3_1
XFILLER_0_79_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_10 _0389_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_21 _0739_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_32 _0912_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_54 _1200_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_65 _1482_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_43 _1038_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_76 _0900_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_87 _1064_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_cap56 _0946_ VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__buf_4
XFILLER_0_38_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2080_ _0739_ _1221_ _1168_ VGND VGND VPWR VPWR _1222_ sky130_fd_sc_hd__a21o_1
XFILLER_0_17_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2982_ _1197_ _0630_ _0631_ _0859_ _0650_ VGND VGND VPWR VPWR _0020_ sky130_fd_sc_hd__o311a_1
XFILLER_0_8_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1933_ net76 VGND VGND VPWR VPWR _0015_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1864_ _0820_ _1007_ _0984_ VGND VGND VPWR VPWR _1008_ sky130_fd_sc_hd__a21o_1
X_1795_ _0939_ _0802_ _0924_ VGND VGND VPWR VPWR _0940_ sky130_fd_sc_hd__and3_4
XFILLER_0_52_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2416_ _0755_ _0832_ _0075_ _0077_ _0694_ VGND VGND VPWR VPWR _0078_ sky130_fd_sc_hd__o311a_1
X_2347_ _1482_ _1483_ _1342_ VGND VGND VPWR VPWR _1484_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2278_ _1367_ _0803_ _0819_ VGND VGND VPWR VPWR _1417_ sky130_fd_sc_hd__and3_1
XFILLER_0_74_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1580_ _0724_ VGND VGND VPWR VPWR _0725_ sky130_fd_sc_hd__buf_4
XFILLER_0_34_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2201_ _1336_ _1338_ _1340_ _1250_ _0843_ VGND VGND VPWR VPWR _1341_ sky130_fd_sc_hd__o221a_1
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2132_ _1193_ VGND VGND VPWR VPWR _1273_ sky130_fd_sc_hd__clkbuf_4
X_2063_ _1204_ _0740_ VGND VGND VPWR VPWR _1205_ sky130_fd_sc_hd__nor2_1
XFILLER_0_88_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2965_ _1367_ _1254_ _0137_ _0957_ VGND VGND VPWR VPWR _0632_ sky130_fd_sc_hd__a211o_1
XFILLER_0_29_397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2896_ _1318_ _0549_ _0551_ _0557_ _1036_ VGND VGND VPWR VPWR _0558_ sky130_fd_sc_hd__o311a_1
XFILLER_0_17_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_507 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1916_ _0984_ VGND VGND VPWR VPWR _1060_ sky130_fd_sc_hd__buf_4
XFILLER_0_44_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1847_ _0937_ _0989_ _0990_ _0967_ _0984_ VGND VGND VPWR VPWR _0991_ sky130_fd_sc_hd__a311o_1
XFILLER_0_8_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1778_ _0922_ VGND VGND VPWR VPWR _0923_ sky130_fd_sc_hd__buf_4
XFILLER_0_12_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_2_3__f_wb_clk_i clknet_0_wb_clk_i VGND VGND VPWR VPWR clknet_2_3__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_94_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_356 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2750_ _1311_ _1213_ _1449_ _0945_ VGND VGND VPWR VPWR _0404_ sky130_fd_sc_hd__a211o_1
XFILLER_0_81_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2681_ _1158_ _0312_ _0313_ _0336_ _0859_ VGND VGND VPWR VPWR _0010_ sky130_fd_sc_hd__o311a_1
X_1701_ net8 net9 _0570_ net10 VGND VGND VPWR VPWR _0846_ sky130_fd_sc_hd__a31o_1
XFILLER_0_53_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1632_ _0776_ VGND VGND VPWR VPWR _0777_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_41_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1563_ _0703_ VGND VGND VPWR VPWR _0706_ sky130_fd_sc_hd__buf_4
XTAP_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3095_ clknet_2_1__leaf_wb_clk_i _0002_ _0030_ VGND VGND VPWR VPWR fsm_inst.done
+ sky130_fd_sc_hd__dfrtp_1
X_2115_ _0836_ VGND VGND VPWR VPWR _1256_ sky130_fd_sc_hd__buf_4
XFILLER_0_89_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2046_ _0784_ _0829_ VGND VGND VPWR VPWR _1188_ sky130_fd_sc_hd__nand2_2
XFILLER_0_49_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2948_ _0834_ _1247_ _1306_ VGND VGND VPWR VPWR _0615_ sky130_fd_sc_hd__or3_1
XFILLER_0_44_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_326 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2879_ _1078_ _1221_ _0959_ _0931_ _0749_ VGND VGND VPWR VPWR _0540_ sky130_fd_sc_hd__a221o_1
XFILLER_0_44_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_112 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2802_ _1199_ _1219_ _0947_ _1172_ _0957_ VGND VGND VPWR VPWR _0457_ sky130_fd_sc_hd__a311o_1
X_2733_ _0383_ _0384_ _0386_ _1342_ _0843_ VGND VGND VPWR VPWR _0387_ sky130_fd_sc_hd__a221o_1
XFILLER_0_42_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2664_ _1190_ _1456_ _1274_ VGND VGND VPWR VPWR _0320_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_41_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2595_ _0667_ _0244_ _0246_ _0248_ _0252_ VGND VGND VPWR VPWR _0253_ sky130_fd_sc_hd__o32a_2
X_1615_ _0759_ VGND VGND VPWR VPWR _0760_ sky130_fd_sc_hd__buf_8
X_1546_ net7 net9 VGND VGND VPWR VPWR _0559_ sky130_fd_sc_hd__and2_1
XFILLER_0_1_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3078_ _0707_ VGND VGND VPWR VPWR _0045_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2029_ _1165_ _1106_ _1166_ _1170_ _0703_ VGND VGND VPWR VPWR _1171_ sky130_fd_sc_hd__o311a_1
XFILLER_0_49_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2380_ _0911_ _0990_ _1516_ VGND VGND VPWR VPWR _1517_ sky130_fd_sc_hd__or3_1
XFILLER_0_36_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3001_ _0663_ VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__buf_1
Xinput6 net80 VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__buf_4
XFILLER_0_78_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2716_ _0873_ _0805_ _0273_ _0370_ _0934_ VGND VGND VPWR VPWR _0371_ sky130_fd_sc_hd__o311a_1
XFILLER_0_14_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2647_ _0741_ _0728_ net54 VGND VGND VPWR VPWR _0303_ sky130_fd_sc_hd__and3_2
XFILLER_0_65_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2578_ _1089_ _1199_ _1019_ _1276_ _1109_ VGND VGND VPWR VPWR _0236_ sky130_fd_sc_hd__a311o_1
XFILLER_0_10_395 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1880_ _1022_ _1023_ _0801_ VGND VGND VPWR VPWR _1024_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_22_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2501_ _1063_ _0733_ _0105_ _0160_ _0950_ VGND VGND VPWR VPWR _0161_ sky130_fd_sc_hd__o311a_1
XFILLER_0_11_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2432_ _0965_ _1275_ _0093_ _1083_ _0914_ VGND VGND VPWR VPWR _0094_ sky130_fd_sc_hd__o221a_1
X_2363_ _1089_ _0713_ _0744_ VGND VGND VPWR VPWR _1500_ sky130_fd_sc_hd__and3_2
X_2294_ _0728_ _1078_ _0996_ VGND VGND VPWR VPWR _1432_ sky130_fd_sc_hd__and3_4
XFILLER_0_59_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_22 _0764_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_11 _0424_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_44 _1072_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_33 _0926_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_66 _1491_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_55 _1202_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_77 _0926_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_284 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_cap57 _0766_ VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__buf_4
XFILLER_0_38_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2981_ _0638_ _0649_ _1197_ VGND VGND VPWR VPWR _0650_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_33_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1932_ net66 _1038_ _1075_ VGND VGND VPWR VPWR _1076_ sky130_fd_sc_hd__and3_1
XFILLER_0_56_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1863_ _0765_ _0760_ VGND VGND VPWR VPWR _1007_ sky130_fd_sc_hd__nor2_4
XFILLER_0_71_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1794_ _0727_ VGND VGND VPWR VPWR _0939_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2415_ _0984_ _1202_ _0076_ VGND VGND VPWR VPWR _0077_ sky130_fd_sc_hd__or3_1
XFILLER_0_58_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2346_ _1160_ _1344_ _1291_ VGND VGND VPWR VPWR _1483_ sky130_fd_sc_hd__a21o_1
X_2277_ _1348_ _0925_ _1380_ _1415_ _1310_ VGND VGND VPWR VPWR _1416_ sky130_fd_sc_hd__o311a_1
Xclkbuf_2_2__f_wb_clk_i clknet_0_wb_clk_i VGND VGND VPWR VPWR clknet_2_2__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_254 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_298 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2200_ _1165_ _0938_ _1141_ _1339_ _1127_ VGND VGND VPWR VPWR _1340_ sky130_fd_sc_hd__o32a_2
X_2131_ _1243_ _1251_ _1258_ _1271_ _0655_ VGND VGND VPWR VPWR _1272_ sky130_fd_sc_hd__o311a_1
XFILLER_0_28_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2062_ _0735_ _0793_ VGND VGND VPWR VPWR _1204_ sky130_fd_sc_hd__nor2_2
XFILLER_0_88_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2964_ _0625_ _0629_ _0655_ VGND VGND VPWR VPWR _0631_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_17_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1915_ _0728_ _0901_ VGND VGND VPWR VPWR _1059_ sky130_fd_sc_hd__nor2_8
XFILLER_0_60_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2895_ _0839_ _0553_ _0556_ _0842_ VGND VGND VPWR VPWR _0557_ sky130_fd_sc_hd__a211o_1
XFILLER_0_56_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1846_ _0740_ _0896_ VGND VGND VPWR VPWR _0990_ sky130_fd_sc_hd__nor2_4
X_1777_ _0799_ VGND VGND VPWR VPWR _0922_ sky130_fd_sc_hd__buf_6
XFILLER_0_69_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2329_ _0772_ _0758_ _0790_ VGND VGND VPWR VPWR _1467_ sky130_fd_sc_hd__and3_2
XFILLER_0_67_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1700_ _0602_ _0623_ VGND VGND VPWR VPWR _0845_ sky130_fd_sc_hd__nand2_1
X_2680_ _0324_ _0335_ _1197_ VGND VGND VPWR VPWR _0336_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_53_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1631_ _0441_ _0679_ VGND VGND VPWR VPWR _0776_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_30_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1562_ _0694_ VGND VGND VPWR VPWR _0703_ sky130_fd_sc_hd__buf_4
XFILLER_0_1_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2114_ _1136_ _1254_ VGND VGND VPWR VPWR _1255_ sky130_fd_sc_hd__nor2_1
XFILLER_0_89_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3094_ clknet_2_0__leaf_wb_clk_i _0001_ _0029_ VGND VGND VPWR VPWR fsm_inst.batch_norm_en
+ sky130_fd_sc_hd__dfrtp_1
X_2045_ _0918_ _0823_ net54 _0864_ VGND VGND VPWR VPWR _1187_ sky130_fd_sc_hd__a31o_2
XFILLER_0_89_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2947_ _1011_ _0787_ _1354_ _1028_ VGND VGND VPWR VPWR _0614_ sky130_fd_sc_hd__a211o_1
XFILLER_0_44_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_338 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2878_ _1040_ _1059_ _0289_ _0538_ _1047_ VGND VGND VPWR VPWR _0539_ sky130_fd_sc_hd__o311a_2
XFILLER_0_13_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1829_ _0972_ VGND VGND VPWR VPWR _0973_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_13_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2801_ _1274_ _1045_ _1094_ _0455_ _0935_ VGND VGND VPWR VPWR _0456_ sky130_fd_sc_hd__o311a_1
XFILLER_0_41_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2732_ _1291_ _0181_ _0186_ _0385_ VGND VGND VPWR VPWR _0386_ sky130_fd_sc_hd__a31o_1
XFILLER_0_26_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2663_ _0755_ _0805_ _1016_ _1330_ VGND VGND VPWR VPWR _0319_ sky130_fd_sc_hd__or4_1
X_2594_ _0915_ _0250_ _0251_ _0842_ VGND VGND VPWR VPWR _0252_ sky130_fd_sc_hd__a31o_1
XFILLER_0_22_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1614_ net3 _0717_ VGND VGND VPWR VPWR _0759_ sky130_fd_sc_hd__and2b_1
XFILLER_0_10_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1545_ _0527_ _0537_ VGND VGND VPWR VPWR _0548_ sky130_fd_sc_hd__nand2_2
XFILLER_0_5_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3077_ _0707_ VGND VGND VPWR VPWR _0044_ sky130_fd_sc_hd__inv_2
XTAP_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2028_ _1167_ _1169_ _0725_ VGND VGND VPWR VPWR _1170_ sky130_fd_sc_hd__a21o_1
XFILLER_0_92_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3000_ weights_inst.data_out\[7\] _0654_ VGND VGND VPWR VPWR _0663_ sky130_fd_sc_hd__and2_1
Xinput7 net82 VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_36_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2715_ _1013_ _0827_ _0929_ _0960_ _0964_ VGND VGND VPWR VPWR _0370_ sky130_fd_sc_hd__a221o_1
X_2646_ _0811_ _0154_ _0173_ VGND VGND VPWR VPWR _0302_ sky130_fd_sc_hd__or3_1
XFILLER_0_77_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2577_ _1259_ _1004_ _1112_ _1151_ _1285_ VGND VGND VPWR VPWR _0235_ sky130_fd_sc_hd__o221a_1
XFILLER_0_10_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3129_ net43 VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__buf_1
XTAP_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_195 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_282 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2500_ _0975_ _0788_ _1059_ _0881_ _0910_ VGND VGND VPWR VPWR _0160_ sky130_fd_sc_hd__a221o_1
X_2431_ _0716_ _0896_ _1052_ VGND VGND VPWR VPWR _0093_ sky130_fd_sc_hd__or3_2
XFILLER_0_11_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2362_ _1345_ _0898_ _0948_ _1498_ _1287_ VGND VGND VPWR VPWR _1499_ sky130_fd_sc_hd__o311a_1
X_2293_ _0985_ _1200_ _1302_ _1430_ _0777_ VGND VGND VPWR VPWR _1431_ sky130_fd_sc_hd__o311a_1
XFILLER_0_79_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_2_1__f_wb_clk_i clknet_0_wb_clk_i VGND VGND VPWR VPWR clknet_2_1__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_74_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_12 _0434_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_23 _0770_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_34 _0965_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_45 _1088_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_56 _1213_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_78 _0948_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_67 _1494_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2629_ _1396_ _0262_ _0269_ _0277_ _0285_ VGND VGND VPWR VPWR _0286_ sky130_fd_sc_hd__o32a_1
XFILLER_0_100_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_cap58 _0452_ VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__buf_4
XFILLER_0_77_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_366 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2980_ _1161_ _0644_ _0648_ VGND VGND VPWR VPWR _0649_ sky130_fd_sc_hd__and3_1
X_1931_ _1039_ _1071_ net75 _0863_ VGND VGND VPWR VPWR _1075_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_33_78 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1862_ _0923_ _0997_ _1002_ _0839_ _1005_ VGND VGND VPWR VPWR _1006_ sky130_fd_sc_hd__o311a_1
XFILLER_0_56_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput10 net64 VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_2
X_1793_ _0918_ _0738_ _0937_ VGND VGND VPWR VPWR _0938_ sky130_fd_sc_hd__and3_2
X_2414_ _0765_ _0784_ _0719_ VGND VGND VPWR VPWR _0076_ sky130_fd_sc_hd__and3_2
X_2345_ _0911_ _0774_ _1467_ VGND VGND VPWR VPWR _1482_ sky130_fd_sc_hd__or3_2
XFILLER_0_74_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2276_ _0917_ _0816_ _1042_ _1264_ VGND VGND VPWR VPWR _1415_ sky130_fd_sc_hd__a211o_1
XFILLER_0_74_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_252 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2130_ _1243_ _1270_ VGND VGND VPWR VPWR _1271_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2061_ _1000_ _0816_ _1202_ _0945_ VGND VGND VPWR VPWR _1203_ sky130_fd_sc_hd__a211o_1
XFILLER_0_88_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2963_ _1396_ _1181_ _0625_ _0629_ VGND VGND VPWR VPWR _0630_ sky130_fd_sc_hd__o211a_1
XFILLER_0_72_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1914_ _1051_ _1057_ _0703_ VGND VGND VPWR VPWR _1058_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_71_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2894_ _1060_ _1422_ _0154_ _0555_ _0914_ VGND VGND VPWR VPWR _0556_ sky130_fd_sc_hd__o311a_1
XFILLER_0_4_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1845_ _0742_ _0831_ VGND VGND VPWR VPWR _0989_ sky130_fd_sc_hd__nand2_8
X_1776_ _0911_ _0912_ _0913_ _0915_ _0920_ VGND VGND VPWR VPWR _0921_ sky130_fd_sc_hd__o311a_1
XFILLER_0_4_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_391 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2328_ _1159_ _1032_ VGND VGND VPWR VPWR _1466_ sky130_fd_sc_hd__and2b_4
X_2259_ _1365_ _1383_ _1397_ VGND VGND VPWR VPWR _1398_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_67_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_58 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1630_ _0767_ _0774_ VGND VGND VPWR VPWR _0775_ sky130_fd_sc_hd__nor2_2
XFILLER_0_22_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1561_ _0685_ VGND VGND VPWR VPWR _0694_ sky130_fd_sc_hd__buf_4
XFILLER_0_1_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2113_ _1123_ _0924_ VGND VGND VPWR VPWR _1254_ sky130_fd_sc_hd__nand2_1
X_3093_ clknet_2_1__leaf_wb_clk_i _0003_ _0028_ VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2044_ _1180_ _0756_ _1182_ _1185_ VGND VGND VPWR VPWR _1186_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_89_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2946_ _1136_ _1031_ _0983_ _0931_ _0956_ VGND VGND VPWR VPWR _0612_ sky130_fd_sc_hd__a221o_1
XFILLER_0_29_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2877_ _1229_ _1399_ _1380_ _1083_ VGND VGND VPWR VPWR _0538_ sky130_fd_sc_hd__a211o_1
XFILLER_0_88_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1828_ _0711_ _0959_ VGND VGND VPWR VPWR _0972_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1759_ _0826_ _0903_ VGND VGND VPWR VPWR _0904_ sky130_fd_sc_hd__or2_1
XFILLER_0_40_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2800_ _1343_ _1020_ _1055_ _0811_ VGND VGND VPWR VPWR _0455_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_41_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2731_ _1199_ _0340_ _0256_ _1211_ VGND VGND VPWR VPWR _0385_ sky130_fd_sc_hd__o211a_1
XFILLER_0_81_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2662_ _0977_ _0316_ _0317_ _1285_ VGND VGND VPWR VPWR _0318_ sky130_fd_sc_hd__o211a_1
XFILLER_0_10_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1613_ _0757_ VGND VGND VPWR VPWR _0758_ sky130_fd_sc_hd__clkbuf_8
X_2593_ _1000_ _0815_ _1266_ _1049_ VGND VGND VPWR VPWR _0251_ sky130_fd_sc_hd__a211o_1
XFILLER_0_10_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1544_ net8 net10 VGND VGND VPWR VPWR _0537_ sky130_fd_sc_hd__or2_2
XFILLER_0_66_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3076_ _0707_ VGND VGND VPWR VPWR _0043_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2027_ _0890_ _1168_ VGND VGND VPWR VPWR _1169_ sky130_fd_sc_hd__nor2_1
XFILLER_0_82_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2929_ _0716_ _0924_ _0959_ VGND VGND VPWR VPWR _0594_ sky130_fd_sc_hd__and3_1
XFILLER_0_33_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_2_0__f_wb_clk_i clknet_0_wb_clk_i VGND VGND VPWR VPWR clknet_2_0__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
Xinput8 net77 VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_78_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2714_ _1403_ _1079_ _0154_ _0368_ _1308_ VGND VGND VPWR VPWR _0369_ sky130_fd_sc_hd__o311a_1
XFILLER_0_2_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2645_ _1124_ _0816_ _1142_ _1281_ VGND VGND VPWR VPWR _0301_ sky130_fd_sc_hd__a211o_1
X_2576_ _1403_ _1174_ _1432_ _0233_ _1308_ VGND VGND VPWR VPWR _0234_ sky130_fd_sc_hd__o311a_1
XFILLER_0_10_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3128_ net43 VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__buf_1
XFILLER_0_96_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3059_ net1 VGND VGND VPWR VPWR _0705_ sky130_fd_sc_hd__buf_4
XFILLER_0_92_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2430_ _0875_ _1189_ _1380_ _0091_ VGND VGND VPWR VPWR _0092_ sky130_fd_sc_hd__o31ai_1
X_2361_ _1335_ _1107_ _1497_ VGND VGND VPWR VPWR _1498_ sky130_fd_sc_hd__nand3_1
X_2292_ _1067_ _1401_ _0754_ VGND VGND VPWR VPWR _1430_ sky130_fd_sc_hd__a21o_1
XFILLER_0_2_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_13 _0449_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_46 _1102_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_35 _0965_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_24 _0787_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_57 _1253_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_68 _0193_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_79 _1041_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2628_ _1164_ _0281_ _0284_ _1039_ VGND VGND VPWR VPWR _0285_ sky130_fd_sc_hd__a31o_1
XFILLER_0_30_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2559_ _1298_ _0208_ _0211_ _0217_ _0861_ VGND VGND VPWR VPWR _0218_ sky130_fd_sc_hd__o311a_1
XFILLER_0_84_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1930_ _0803_ _1072_ _1053_ _1073_ _1036_ VGND VGND VPWR VPWR _1074_ sky130_fd_sc_hd__a221o_1
XFILLER_0_29_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1861_ _0824_ _0807_ _1004_ _0836_ VGND VGND VPWR VPWR _1005_ sky130_fd_sc_hd__a211o_1
XFILLER_0_56_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput11 net84 VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__clkbuf_1
X_1792_ _0771_ _0886_ VGND VGND VPWR VPWR _0937_ sky130_fd_sc_hd__nand2_4
XFILLER_0_12_437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2413_ _0728_ _1181_ VGND VGND VPWR VPWR _0075_ sky130_fd_sc_hd__nor2_4
XFILLER_0_20_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2344_ _1347_ _1088_ _1054_ VGND VGND VPWR VPWR _1481_ sky130_fd_sc_hd__o21ai_1
X_2275_ _1298_ _1404_ _1406_ _1413_ _1396_ VGND VGND VPWR VPWR _1414_ sky130_fd_sc_hd__o311a_1
XFILLER_0_74_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2060_ _0768_ _0989_ VGND VGND VPWR VPWR _1202_ sky130_fd_sc_hd__and2_4
XFILLER_0_88_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2962_ _1250_ _0583_ _0626_ _0628_ _1164_ VGND VGND VPWR VPWR _0629_ sky130_fd_sc_hd__a311o_1
XFILLER_0_56_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1913_ _1054_ _1055_ _1056_ VGND VGND VPWR VPWR _1057_ sky130_fd_sc_hd__a21o_1
XFILLER_0_44_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2893_ _0723_ _0890_ _1168_ _0554_ VGND VGND VPWR VPWR _0555_ sky130_fd_sc_hd__or4_1
XFILLER_0_71_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1844_ _0758_ _0937_ _0947_ VGND VGND VPWR VPWR _0988_ sky130_fd_sc_hd__and3_4
XFILLER_0_4_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1775_ _0917_ _0919_ _0875_ VGND VGND VPWR VPWR _0920_ sky130_fd_sc_hd__a21o_1
XFILLER_0_4_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2327_ _0985_ _1407_ _1462_ _1464_ _0838_ VGND VGND VPWR VPWR _1465_ sky130_fd_sc_hd__o311a_1
X_2258_ _1298_ _1386_ _1388_ _1395_ _1396_ VGND VGND VPWR VPWR _1397_ sky130_fd_sc_hd__o311a_1
XFILLER_0_33_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2189_ _0918_ _0903_ VGND VGND VPWR VPWR _1329_ sky130_fd_sc_hd__nand2_2
XFILLER_0_67_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1560_ _0441_ _0679_ VGND VGND VPWR VPWR _0685_ sky130_fd_sc_hd__xor2_4
XFILLER_0_22_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2112_ _0799_ _1252_ VGND VGND VPWR VPWR _1253_ sky130_fd_sc_hd__or2_4
X_3092_ net1 VGND VGND VPWR VPWR _0058_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2043_ _0835_ _0733_ _1183_ _1184_ VGND VGND VPWR VPWR _1185_ sky130_fd_sc_hd__or4_1
XFILLER_0_9_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2945_ _0875_ _1206_ _1130_ _0610_ _0934_ VGND VGND VPWR VPWR _0611_ sky130_fd_sc_hd__o311a_1
X_2876_ _1109_ _1432_ _0467_ _0535_ _0978_ VGND VGND VPWR VPWR _0536_ sky130_fd_sc_hd__o311a_1
X_1827_ _0797_ VGND VGND VPWR VPWR _0971_ sky130_fd_sc_hd__buf_4
XFILLER_0_4_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1758_ _0741_ _0742_ _0718_ VGND VGND VPWR VPWR _0903_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_40_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1689_ _0833_ VGND VGND VPWR VPWR _0834_ sky130_fd_sc_hd__clkbuf_4
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_392 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2730_ _1391_ _0744_ _1147_ _0915_ VGND VGND VPWR VPWR _0384_ sky130_fd_sc_hd__o31a_1
XFILLER_0_81_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2661_ _1073_ _1379_ _1137_ _0801_ VGND VGND VPWR VPWR _0317_ sky130_fd_sc_hd__a211o_1
X_1612_ _0715_ VGND VGND VPWR VPWR _0757_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_22_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2592_ _1065_ _0249_ _1063_ VGND VGND VPWR VPWR _0250_ sky130_fd_sc_hd__a21o_1
XFILLER_0_10_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1543_ net8 net10 VGND VGND VPWR VPWR _0527_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_395 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3075_ _0707_ VGND VGND VPWR VPWR _0042_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2026_ net58 _0976_ VGND VGND VPWR VPWR _1168_ sky130_fd_sc_hd__nor2_2
XFILLER_0_82_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2928_ _0964_ _1276_ _0590_ _0592_ _0777_ VGND VGND VPWR VPWR _0593_ sky130_fd_sc_hd__o311a_1
XFILLER_0_72_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2859_ _1298_ _0510_ _0512_ _0518_ VGND VGND VPWR VPWR _0519_ sky130_fd_sc_hd__a31o_1
XFILLER_0_32_115 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_270 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput9 net68 VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__buf_4
XFILLER_0_36_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2713_ _1367_ _0824_ _0807_ _1020_ _1040_ VGND VGND VPWR VPWR _0368_ sky130_fd_sc_hd__a221o_1
X_2644_ _1322_ _0286_ _0300_ _1242_ VGND VGND VPWR VPWR _0009_ sky130_fd_sc_hd__o211a_1
XFILLER_0_42_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2575_ _0936_ _1162_ _1288_ VGND VGND VPWR VPWR _0233_ sky130_fd_sc_hd__or3_1
XFILLER_0_2_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3127_ net43 VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__buf_1
XFILLER_0_89_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3058_ _0695_ _0700_ _0704_ VGND VGND VPWR VPWR fsm_inst.next_state\[2\] sky130_fd_sc_hd__o21ai_1
XFILLER_0_65_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2009_ _0716_ _0924_ _0851_ VGND VGND VPWR VPWR _1152_ sky130_fd_sc_hd__and3_2
XFILLER_0_92_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_251 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2360_ _0769_ _1073_ VGND VGND VPWR VPWR _1497_ sky130_fd_sc_hd__or2_2
X_2291_ _1158_ _1398_ _1429_ _1242_ VGND VGND VPWR VPWR _0024_ sky130_fd_sc_hd__o211a_1
XFILLER_0_63_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_14 _0467_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_47 _1103_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_25 _0798_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_36 _0990_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_69 _0733_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_58 _1307_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2627_ _0915_ _0282_ _0283_ VGND VGND VPWR VPWR _0284_ sky130_fd_sc_hd__or3b_1
X_2558_ _1310_ _0212_ _0213_ _0216_ _1318_ VGND VGND VPWR VPWR _0217_ sky130_fd_sc_hd__a311o_1
X_2489_ _0779_ _0144_ _0145_ _0148_ _0667_ VGND VGND VPWR VPWR _0149_ sky130_fd_sc_hd__a311o_1
XFILLER_0_97_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1860_ _1003_ _0785_ VGND VGND VPWR VPWR _1004_ sky130_fd_sc_hd__and2_1
XFILLER_0_71_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1791_ _0910_ VGND VGND VPWR VPWR _0936_ sky130_fd_sc_hd__buf_4
Xinput12 wbs_cyc_i VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2412_ _1287_ _0069_ _0070_ _0073_ VGND VGND VPWR VPWR _0074_ sky130_fd_sc_hd__a31o_1
X_2343_ _1480_ VGND VGND VPWR VPWR _0025_ sky130_fd_sc_hd__clkbuf_1
X_2274_ _0779_ _1408_ _1409_ _1412_ _0667_ VGND VGND VPWR VPWR _1413_ sky130_fd_sc_hd__a311o_1
XFILLER_0_79_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1989_ _0944_ _1066_ _1129_ _1131_ _0777_ VGND VGND VPWR VPWR _1132_ sky130_fd_sc_hd__o311a_1
XFILLER_0_43_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2961_ _0811_ _0627_ _0585_ _0839_ VGND VGND VPWR VPWR _0628_ sky130_fd_sc_hd__o211a_1
XFILLER_0_56_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1912_ _0724_ VGND VGND VPWR VPWR _1056_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_8_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_327 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2892_ _0772_ _0712_ _0826_ VGND VGND VPWR VPWR _0554_ sky130_fd_sc_hd__a21oi_1
X_1843_ _0898_ _0899_ _0936_ VGND VGND VPWR VPWR _0987_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_25_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1774_ _0881_ _0819_ _0918_ VGND VGND VPWR VPWR _0919_ sky130_fd_sc_hd__a21o_2
XFILLER_0_52_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2326_ _1123_ _1106_ _1463_ _0799_ VGND VGND VPWR VPWR _1464_ sky130_fd_sc_hd__a211o_1
XTAP_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2257_ _1036_ VGND VGND VPWR VPWR _1396_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_26_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2188_ _1261_ _1202_ _1323_ _1327_ _1178_ VGND VGND VPWR VPWR _1328_ sky130_fd_sc_hd__o311a_1
XFILLER_0_79_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1 wbs_dat_i[0] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__dlygate4sd3_1
X_3091_ _0709_ VGND VGND VPWR VPWR _0057_ sky130_fd_sc_hd__inv_2
X_2111_ _0826_ _1064_ VGND VGND VPWR VPWR _1252_ sky130_fd_sc_hd__nor2_2
X_2042_ _0745_ _0887_ _0959_ VGND VGND VPWR VPWR _1184_ sky130_fd_sc_hd__and3_2
XFILLER_0_55_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2944_ _1013_ _1106_ _0303_ _0944_ VGND VGND VPWR VPWR _0610_ sky130_fd_sc_hd__a211o_1
XFILLER_0_72_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2875_ _0724_ _0747_ _1277_ VGND VGND VPWR VPWR _0535_ sky130_fd_sc_hd__or3_1
XFILLER_0_72_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1826_ _0926_ VGND VGND VPWR VPWR _0970_ sky130_fd_sc_hd__buf_4
XFILLER_0_4_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1757_ _0756_ _0768_ _0719_ _0813_ net58 VGND VGND VPWR VPWR _0902_ sky130_fd_sc_hd__a32o_1
XFILLER_0_96_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1688_ _0473_ _0505_ VGND VGND VPWR VPWR _0833_ sky130_fd_sc_hd__xor2_2
XFILLER_0_96_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2309_ _1445_ _1446_ _0915_ VGND VGND VPWR VPWR _1447_ sky130_fd_sc_hd__a21oi_1
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_474 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2660_ _1261_ _1329_ VGND VGND VPWR VPWR _0316_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1611_ _0711_ _0737_ VGND VGND VPWR VPWR _0756_ sky130_fd_sc_hd__xnor2_4
X_2591_ _0769_ _0989_ _1325_ _0854_ VGND VGND VPWR VPWR _0249_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1542_ _0441_ _0473_ _0505_ VGND VGND VPWR VPWR _0516_ sky130_fd_sc_hd__and3_4
XFILLER_0_10_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3074_ _0707_ VGND VGND VPWR VPWR _0041_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2025_ _0785_ _0870_ VGND VGND VPWR VPWR _1167_ sky130_fd_sc_hd__nand2_4
XFILLER_0_89_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_135 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2927_ _0825_ _1077_ _0137_ _0749_ VGND VGND VPWR VPWR _0592_ sky130_fd_sc_hd__a211o_1
XFILLER_0_93_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2858_ _0907_ _0514_ _0517_ _0860_ VGND VGND VPWR VPWR _0518_ sky130_fd_sc_hd__a31o_1
XFILLER_0_5_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1809_ _0843_ _0921_ _0933_ _0953_ _0863_ VGND VGND VPWR VPWR _0954_ sky130_fd_sc_hd__o311a_1
X_2789_ _1391_ _1078_ VGND VGND VPWR VPWR _0444_ sky130_fd_sc_hd__nor2_1
XFILLER_0_40_171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_282 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2712_ _0787_ _1259_ _1044_ _0366_ _0779_ VGND VGND VPWR VPWR _0367_ sky130_fd_sc_hd__o311a_1
XFILLER_0_42_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2643_ _0298_ _0299_ _1322_ VGND VGND VPWR VPWR _0300_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_2_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2574_ _0220_ _0231_ VGND VGND VPWR VPWR _0232_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_97_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3126_ net43 VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__buf_1
XTAP_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3057_ fsm_inst.current_state\[1\] _0701_ _0702_ _0002_ VGND VGND VPWR VPWR _0704_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_89_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2008_ _0820_ _0823_ net54 _0799_ VGND VGND VPWR VPWR _1151_ sky130_fd_sc_hd__a31o_2
XFILLER_0_65_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2290_ _1414_ _1428_ _1197_ VGND VGND VPWR VPWR _1429_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_47_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_37 _1001_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_26 _0840_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_15 _0560_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_48 _1103_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_59 _1354_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2626_ _0786_ _0965_ _1399_ _0807_ _0836_ VGND VGND VPWR VPWR _0283_ sky130_fd_sc_hd__a221o_1
XFILLER_0_30_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2557_ _0945_ _1175_ _0214_ _0215_ _0978_ VGND VGND VPWR VPWR _0216_ sky130_fd_sc_hd__o311a_1
XFILLER_0_56_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2488_ _1056_ _0980_ _0146_ _0147_ _0963_ VGND VGND VPWR VPWR _0148_ sky130_fd_sc_hd__o311a_1
XFILLER_0_97_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3109_ clknet_2_2__leaf_wb_clk_i _0027_ _0044_ VGND VGND VPWR VPWR weights_inst.data_out\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput13 net60 VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__buf_1
X_1790_ _0934_ VGND VGND VPWR VPWR _0935_ sky130_fd_sc_hd__buf_4
XFILLER_0_24_222 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2411_ _0934_ _0071_ _0072_ _0661_ VGND VGND VPWR VPWR _0073_ sky130_fd_sc_hd__a31o_1
X_2342_ _1479_ _0859_ VGND VGND VPWR VPWR _1480_ sky130_fd_sc_hd__and2b_1
X_2273_ _0945_ _1119_ _1410_ _1411_ _0963_ VGND VGND VPWR VPWR _1412_ sky130_fd_sc_hd__o311a_1
XFILLER_0_74_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1988_ _0749_ _1027_ _1130_ VGND VGND VPWR VPWR _1131_ sky130_fd_sc_hd__or3_1
XFILLER_0_43_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2609_ _0939_ _0738_ _0924_ VGND VGND VPWR VPWR _0266_ sky130_fd_sc_hd__and3_2
XFILLER_0_11_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2960_ _0771_ _1146_ _0744_ VGND VGND VPWR VPWR _0627_ sky130_fd_sc_hd__a21oi_1
XTAP_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2891_ _1089_ _1083_ _0770_ _0552_ _1124_ VGND VGND VPWR VPWR _0553_ sky130_fd_sc_hd__a32o_1
X_1911_ _0737_ _0877_ VGND VGND VPWR VPWR _1055_ sky130_fd_sc_hd__nand2_4
XFILLER_0_84_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1842_ _0916_ _0815_ _0983_ _0931_ _0985_ VGND VGND VPWR VPWR _0986_ sky130_fd_sc_hd__a221o_1
XFILLER_0_44_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1773_ _0826_ VGND VGND VPWR VPWR _0918_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_69_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2325_ _0791_ _0805_ VGND VGND VPWR VPWR _1463_ sky130_fd_sc_hd__nor2_1
XTAP_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2256_ _1285_ _1389_ _1390_ _1394_ _1318_ VGND VGND VPWR VPWR _1395_ sky130_fd_sc_hd__a311o_1
XFILLER_0_79_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2187_ _1049_ _1324_ _1326_ VGND VGND VPWR VPWR _1327_ sky130_fd_sc_hd__or3_1
XFILLER_0_48_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2 fsm_inst.next_state\[0\] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__dlygate4sd3_1
X_3090_ _0709_ VGND VGND VPWR VPWR _0056_ sky130_fd_sc_hd__inv_2
X_2110_ _1244_ _1246_ _1248_ _1249_ _1250_ VGND VGND VPWR VPWR _1251_ sky130_fd_sc_hd__o221a_1
X_2041_ _0772_ _1015_ VGND VGND VPWR VPWR _1183_ sky130_fd_sc_hd__nor2_4
XFILLER_0_55_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2943_ _0607_ _0608_ _0782_ VGND VGND VPWR VPWR _0609_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_72_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2874_ _1322_ _0520_ _0534_ _1242_ VGND VGND VPWR VPWR _0016_ sky130_fd_sc_hd__o211a_1
XFILLER_0_72_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1825_ _0957_ _0960_ _0962_ _0963_ _0968_ VGND VGND VPWR VPWR _0969_ sky130_fd_sc_hd__o311a_1
X_1756_ _0828_ _0765_ VGND VGND VPWR VPWR _0901_ sky130_fd_sc_hd__nor2_4
XFILLER_0_4_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1687_ _0745_ _0732_ _0829_ _0831_ VGND VGND VPWR VPWR _0832_ sky130_fd_sc_hd__and4_2
XFILLER_0_96_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2308_ _1003_ _0878_ _1013_ _1294_ _0922_ VGND VGND VPWR VPWR _1446_ sky130_fd_sc_hd__a311o_1
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2239_ _1077_ VGND VGND VPWR VPWR _1379_ sky130_fd_sc_hd__buf_4
XFILLER_0_95_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1610_ _0754_ VGND VGND VPWR VPWR _0755_ sky130_fd_sc_hd__buf_6
X_2590_ _1165_ _1229_ _1072_ _0247_ _0839_ VGND VGND VPWR VPWR _0248_ sky130_fd_sc_hd__o311a_1
X_1541_ _0484_ _0495_ VGND VGND VPWR VPWR _0505_ sky130_fd_sc_hd__and2_2
XFILLER_0_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3073_ _0707_ VGND VGND VPWR VPWR _0040_ sky130_fd_sc_hd__inv_2
X_2024_ _1003_ _0769_ VGND VGND VPWR VPWR _1166_ sky130_fd_sc_hd__nor2_2
XFILLER_0_82_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2926_ _0926_ _0713_ _0999_ VGND VGND VPWR VPWR _0590_ sky130_fd_sc_hd__and3_2
XFILLER_0_72_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2857_ _0936_ _0390_ _0186_ _0515_ _0934_ VGND VGND VPWR VPWR _0517_ sky130_fd_sc_hd__a311o_1
XFILLER_0_17_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1808_ _0935_ _0943_ _0951_ _0952_ VGND VGND VPWR VPWR _0953_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_13_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2788_ _0345_ _0724_ _1098_ VGND VGND VPWR VPWR _0443_ sky130_fd_sc_hd__or3b_1
XFILLER_0_60_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1739_ _0875_ _0876_ _0879_ _0883_ VGND VGND VPWR VPWR _0884_ sky130_fd_sc_hd__a31o_1
XFILLER_0_40_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2711_ _1125_ _1334_ _1335_ VGND VGND VPWR VPWR _0366_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_54_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2642_ _0871_ _1065_ _0655_ VGND VGND VPWR VPWR _0299_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_2_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2573_ _0706_ _0223_ _0225_ _0230_ VGND VGND VPWR VPWR _0231_ sky130_fd_sc_hd__o31a_2
XFILLER_0_77_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3125_ net43 VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__buf_1
XFILLER_0_96_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3056_ fsm_inst.current_state\[1\] fsm_inst.current_state\[0\] fsm_inst.current_state\[2\]
+ VGND VGND VPWR VPWR _0702_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_89_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2007_ _0740_ _0831_ _0818_ VGND VGND VPWR VPWR _1150_ sky130_fd_sc_hd__and3_2
XFILLER_0_65_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2909_ _1036_ _0075_ VGND VGND VPWR VPWR _0573_ sky130_fd_sc_hd__nor2_1
XFILLER_0_18_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_38 _1034_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_16 _0608_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_27 _0878_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_49 _1154_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2625_ _1255_ _1049_ _0722_ VGND VGND VPWR VPWR _0282_ sky130_fd_sc_hd__and3b_1
XFILLER_0_88_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2556_ _0724_ _0832_ _1214_ VGND VGND VPWR VPWR _0215_ sky130_fd_sc_hd__or3b_4
X_2487_ _1124_ _1136_ _1078_ _0806_ _1028_ VGND VGND VPWR VPWR _0147_ sky130_fd_sc_hd__a221o_1
XFILLER_0_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3108_ clknet_2_3__leaf_wb_clk_i _0026_ _0043_ VGND VGND VPWR VPWR weights_inst.data_out\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3039_ fsm_inst.current_state\[1\] fsm_inst.current_state\[0\] fsm_inst.current_state\[2\]
+ VGND VGND VPWR VPWR _0687_ sky130_fd_sc_hd__and3_1
XFILLER_0_65_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput14 net62 VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__buf_1
XFILLER_0_24_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2410_ _1089_ _0970_ _0893_ _0750_ VGND VGND VPWR VPWR _0072_ sky130_fd_sc_hd__a211o_1
X_2341_ _1442_ _1444_ _1461_ _1478_ _0863_ _0645_ VGND VGND VPWR VPWR _1479_ sky130_fd_sc_hd__mux4_1
X_2272_ _1011_ _1097_ _1301_ _0750_ VGND VGND VPWR VPWR _1411_ sky130_fd_sc_hd__a211o_1
XFILLER_0_79_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1987_ _0794_ _0727_ _0853_ VGND VGND VPWR VPWR _1130_ sky130_fd_sc_hd__and3_2
XFILLER_0_55_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2608_ _1256_ _1453_ _0264_ _0839_ VGND VGND VPWR VPWR _0265_ sky130_fd_sc_hd__a31o_1
XFILLER_0_30_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2539_ _1348_ _1174_ VGND VGND VPWR VPWR _0198_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2890_ _0724_ _0899_ _1219_ VGND VGND VPWR VPWR _0552_ sky130_fd_sc_hd__o21ai_1
X_1910_ _0802_ _1053_ VGND VGND VPWR VPWR _1054_ sky130_fd_sc_hd__nand2_2
XTAP_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1841_ _0984_ VGND VGND VPWR VPWR _0985_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_44_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1772_ _0916_ VGND VGND VPWR VPWR _0917_ sky130_fd_sc_hd__buf_4
XFILLER_0_8_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2324_ _0854_ _1325_ _1041_ VGND VGND VPWR VPWR _1462_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_85_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2255_ _1175_ _1225_ _1393_ _0963_ VGND VGND VPWR VPWR _1394_ sky130_fd_sc_hd__o211a_1
X_2186_ _0854_ _1325_ _0975_ VGND VGND VPWR VPWR _1326_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_79_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_395 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3 wbs_dat_i[1] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__dlygate4sd3_1
X_2040_ _0770_ _1181_ VGND VGND VPWR VPWR _1182_ sky130_fd_sc_hd__nor2_2
XFILLER_0_69_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2942_ _0910_ _0948_ _0913_ VGND VGND VPWR VPWR _0608_ sky130_fd_sc_hd__or3_4
XFILLER_0_84_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2873_ _0655_ _0526_ _0532_ _0533_ _0849_ VGND VGND VPWR VPWR _0534_ sky130_fd_sc_hd__a311o_1
X_1824_ _0964_ _0966_ _0967_ VGND VGND VPWR VPWR _0968_ sky130_fd_sc_hd__or3_1
X_1755_ _0723_ _0899_ VGND VGND VPWR VPWR _0900_ sky130_fd_sc_hd__or2_4
XFILLER_0_20_61 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1686_ _0830_ VGND VGND VPWR VPWR _0831_ sky130_fd_sc_hd__buf_4
XFILLER_0_40_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2307_ _0835_ _1249_ _1050_ _1410_ VGND VGND VPWR VPWR _1445_ sky130_fd_sc_hd__or4_1
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2238_ _1243_ _1369_ _1371_ _1377_ VGND VGND VPWR VPWR _1378_ sky130_fd_sc_hd__o31a_1
XFILLER_0_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2169_ _1115_ VGND VGND VPWR VPWR _1310_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_67_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1540_ net6 net8 VGND VGND VPWR VPWR _0495_ sky130_fd_sc_hd__or2_1
XFILLER_0_22_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3072_ _0707_ VGND VGND VPWR VPWR _0039_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2023_ _1049_ VGND VGND VPWR VPWR _1165_ sky130_fd_sc_hd__buf_4
XFILLER_0_9_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2925_ _0907_ _0578_ _0582_ _0588_ VGND VGND VPWR VPWR _0589_ sky130_fd_sc_hd__a31o_1
XFILLER_0_45_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2856_ _1060_ _0815_ _1118_ VGND VGND VPWR VPWR _0515_ sky130_fd_sc_hd__nor3_1
XFILLER_0_45_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1807_ _0842_ VGND VGND VPWR VPWR _0952_ sky130_fd_sc_hd__buf_4
XFILLER_0_31_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2787_ _0075_ _0158_ _0440_ _0782_ VGND VGND VPWR VPWR _0442_ sky130_fd_sc_hd__o211a_1
XFILLER_0_13_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1738_ _0864_ _0823_ _0880_ _0882_ VGND VGND VPWR VPWR _0883_ sky130_fd_sc_hd__and4_1
XFILLER_0_40_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1669_ _0768_ _0813_ VGND VGND VPWR VPWR _0814_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2710_ _0645_ _0355_ _0357_ _0364_ _0673_ VGND VGND VPWR VPWR _0365_ sky130_fd_sc_hd__o311a_1
XFILLER_0_42_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2641_ _0673_ _0288_ _0291_ _0297_ _1161_ VGND VGND VPWR VPWR _0298_ sky130_fd_sc_hd__o311a_2
XFILLER_0_2_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2572_ _1193_ _0226_ _0227_ _1178_ _0229_ VGND VGND VPWR VPWR _0230_ sky130_fd_sc_hd__a311o_1
XFILLER_0_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3055_ net13 _0690_ fsm_inst.current_state\[0\] VGND VGND VPWR VPWR _0701_ sky130_fd_sc_hd__a21oi_1
X_2006_ _1031_ _0868_ _1147_ _1148_ _0836_ VGND VGND VPWR VPWR _1149_ sky130_fd_sc_hd__o32a_1
XFILLER_0_77_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2908_ _1318_ _0565_ _0571_ VGND VGND VPWR VPWR _0572_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_73_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2839_ _1055_ _1359_ _0752_ VGND VGND VPWR VPWR _0497_ sky130_fd_sc_hd__a21o_1
XFILLER_0_5_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_438 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_26 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_28 _0888_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_17 _0617_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_39 _1038_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2624_ _0278_ _0279_ _0280_ _1278_ VGND VGND VPWR VPWR _0281_ sky130_fd_sc_hd__a211o_2
XFILLER_0_100_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2555_ _1106_ _1254_ VGND VGND VPWR VPWR _0214_ sky130_fd_sc_hd__and2_1
X_2486_ _0881_ _0939_ _0797_ VGND VGND VPWR VPWR _0146_ sky130_fd_sc_hd__and3_2
X_3107_ clknet_2_0__leaf_wb_clk_i _0025_ _0042_ VGND VGND VPWR VPWR weights_inst.data_out\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_3038_ _0686_ VGND VGND VPWR VPWR _0001_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput15 wbs_dat_i[2] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__buf_1
XFILLER_0_52_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2340_ _0842_ _1465_ _1469_ _1473_ _1477_ VGND VGND VPWR VPWR _1478_ sky130_fd_sc_hd__o32a_1
X_2271_ _1015_ _0961_ VGND VGND VPWR VPWR _1410_ sky130_fd_sc_hd__nor2_4
XFILLER_0_87_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1986_ _0939_ _0797_ _0927_ VGND VGND VPWR VPWR _1129_ sky130_fd_sc_hd__and3_2
XFILLER_0_55_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2607_ _1206_ _1025_ VGND VGND VPWR VPWR _0264_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2538_ _1348_ _0720_ _1249_ _0196_ _1287_ VGND VGND VPWR VPWR _0197_ sky130_fd_sc_hd__o311a_1
X_2469_ _0918_ _0896_ VGND VGND VPWR VPWR _0130_ sky130_fd_sc_hd__nor2_1
XFILLER_0_97_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1840_ _0833_ VGND VGND VPWR VPWR _0984_ sky130_fd_sc_hd__buf_4
XFILLER_0_25_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1771_ _0790_ VGND VGND VPWR VPWR _0916_ sky130_fd_sc_hd__buf_4
XFILLER_0_69_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2323_ _1447_ _1452_ _1460_ VGND VGND VPWR VPWR _1461_ sky130_fd_sc_hd__o21ai_1
XTAP_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2254_ _1020_ _1392_ _1083_ VGND VGND VPWR VPWR _1393_ sky130_fd_sc_hd__a21o_1
XFILLER_0_79_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2185_ _0735_ _0719_ _0737_ VGND VGND VPWR VPWR _1325_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_79_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_382 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1969_ _0826_ _0829_ _0831_ VGND VGND VPWR VPWR _1112_ sky130_fd_sc_hd__and3_2
XFILLER_0_98_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4 fsm_inst.next_state\[1\] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2941_ _0264_ _0093_ _0755_ VGND VGND VPWR VPWR _0607_ sky130_fd_sc_hd__a21o_1
XFILLER_0_29_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_135 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_422 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_466 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2872_ _1124_ _0880_ _1532_ _1039_ VGND VGND VPWR VPWR _0533_ sky130_fd_sc_hd__o211a_1
XFILLER_0_72_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1823_ _0784_ _0719_ _0790_ VGND VGND VPWR VPWR _0967_ sky130_fd_sc_hd__and3_1
X_1754_ _0772_ _0768_ VGND VGND VPWR VPWR _0899_ sky130_fd_sc_hd__nor2_2
XFILLER_0_13_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1685_ _0717_ _0708_ VGND VGND VPWR VPWR _0830_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2306_ _1089_ _1343_ _0929_ _1443_ VGND VGND VPWR VPWR _1444_ sky130_fd_sc_hd__a31o_1
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2237_ _0783_ _1372_ _1373_ _1376_ VGND VGND VPWR VPWR _1377_ sky130_fd_sc_hd__a31o_2
XFILLER_0_24_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2168_ _1281_ _0988_ _1305_ _1307_ _1308_ VGND VGND VPWR VPWR _1309_ sky130_fd_sc_hd__o311a_1
XFILLER_0_95_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2099_ _1197_ _1240_ VGND VGND VPWR VPWR _1241_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xkws_wrapper_59 VGND VGND VPWR VPWR kws_wrapper_59/HI wbs_dat_o[31] sky130_fd_sc_hd__conb_1
XFILLER_0_41_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3071_ _0707_ VGND VGND VPWR VPWR _0038_ sky130_fd_sc_hd__inv_2
X_2022_ _0993_ VGND VGND VPWR VPWR _1164_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2924_ _0584_ _0587_ _0841_ VGND VGND VPWR VPWR _0588_ sky130_fd_sc_hd__o21a_1
XFILLER_0_57_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2855_ _1056_ _0871_ _1055_ _0513_ _0694_ VGND VGND VPWR VPWR _0514_ sky130_fd_sc_hd__a311o_1
XFILLER_0_33_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1806_ _0945_ net56 _0882_ _0949_ _0950_ VGND VGND VPWR VPWR _0951_ sky130_fd_sc_hd__a221o_1
XFILLER_0_60_439 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2786_ _0878_ _1173_ _1466_ _0922_ VGND VGND VPWR VPWR _0440_ sky130_fd_sc_hd__a211o_1
X_1737_ _0881_ _0716_ VGND VGND VPWR VPWR _0882_ sky130_fd_sc_hd__nand2_2
XFILLER_0_40_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1668_ _0812_ VGND VGND VPWR VPWR _0813_ sky130_fd_sc_hd__clkbuf_8
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1599_ _0740_ _0743_ VGND VGND VPWR VPWR _0744_ sky130_fd_sc_hd__nor2_8
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2640_ _1342_ _0294_ _0296_ _0952_ VGND VGND VPWR VPWR _0297_ sky130_fd_sc_hd__a211o_1
XFILLER_0_2_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2571_ _1063_ _1141_ _1302_ _0228_ _0661_ VGND VGND VPWR VPWR _0229_ sky130_fd_sc_hd__o311a_1
XFILLER_0_2_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3123_ clknet_2_3__leaf_wb_clk_i _0020_ _0058_ VGND VGND VPWR VPWR weights_inst.data_out\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_3054_ _0696_ _0690_ VGND VGND VPWR VPWR _0700_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2005_ _1013_ _1106_ _0925_ VGND VGND VPWR VPWR _1148_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_9_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2907_ _0778_ _0566_ _0567_ _0569_ _0841_ VGND VGND VPWR VPWR _0571_ sky130_fd_sc_hd__a311o_1
XFILLER_0_91_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2838_ _1206_ _0172_ _1457_ _1281_ VGND VGND VPWR VPWR _0496_ sky130_fd_sc_hd__a211o_1
XFILLER_0_13_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2769_ _0764_ _0389_ _0964_ VGND VGND VPWR VPWR _0423_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_13_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_18 _0645_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_29 _0888_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2623_ _1261_ _0278_ VGND VGND VPWR VPWR _0280_ sky130_fd_sc_hd__nor2_1
X_2554_ _0725_ _0938_ _0154_ VGND VGND VPWR VPWR _0213_ sky130_fd_sc_hd__or3_1
X_2485_ _1311_ _1219_ _0947_ _1166_ _1180_ VGND VGND VPWR VPWR _0145_ sky130_fd_sc_hd__a311o_1
X_3106_ clknet_2_2__leaf_wb_clk_i _0024_ _0041_ VGND VGND VPWR VPWR weights_inst.data_out\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3037_ fsm_inst.current_state\[0\] fsm_inst.current_state\[2\] fsm_inst.current_state\[1\]
+ VGND VGND VPWR VPWR _0686_ sky130_fd_sc_hd__and3b_1
XFILLER_0_93_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_391 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_247 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput16 wbs_dat_i[3] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__buf_1
XFILLER_0_37_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_59 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2270_ _1073_ _1379_ _1180_ _1066_ VGND VGND VPWR VPWR _1409_ sky130_fd_sc_hd__a211o_1
XFILLER_0_59_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1985_ _0999_ _0916_ _1084_ _1127_ _0750_ VGND VGND VPWR VPWR _1128_ sky130_fd_sc_hd__a311o_1
XFILLER_0_99_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2606_ _1343_ _0195_ _1001_ _1124_ _1291_ VGND VGND VPWR VPWR _0263_ sky130_fd_sc_hd__o221a_1
XFILLER_0_101_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2537_ _1211_ _0195_ _1407_ VGND VGND VPWR VPWR _0196_ sky130_fd_sc_hd__or3_1
X_2468_ _0739_ _0817_ _1220_ _0128_ VGND VGND VPWR VPWR _0129_ sky130_fd_sc_hd__a31o_1
XFILLER_0_54_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2399_ _1274_ _1042_ _1129_ _0060_ _1278_ VGND VGND VPWR VPWR _0061_ sky130_fd_sc_hd__o311a_1
XFILLER_0_97_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_383 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1770_ _0914_ VGND VGND VPWR VPWR _0915_ sky130_fd_sc_hd__buf_4
XFILLER_0_40_504 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2322_ _0934_ _1455_ _1459_ _0661_ VGND VGND VPWR VPWR _1460_ sky130_fd_sc_hd__a211o_1
XFILLER_0_20_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2253_ _0726_ _1391_ _1031_ VGND VGND VPWR VPWR _1392_ sky130_fd_sc_hd__or3_4
X_2184_ _0768_ _0886_ VGND VGND VPWR VPWR _1324_ sky130_fd_sc_hd__nor2_4
XFILLER_0_79_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_0_wb_clk_i wb_clk_i VGND VGND VPWR VPWR clknet_0_wb_clk_i sky130_fd_sc_hd__clkbuf_16
XFILLER_0_94_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_394 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1968_ _0743_ _1110_ VGND VGND VPWR VPWR _1111_ sky130_fd_sc_hd__nor2_2
XFILLER_0_16_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1899_ _1032_ VGND VGND VPWR VPWR _1043_ sky130_fd_sc_hd__buf_4
XFILLER_0_3_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold5 wbs_adr_i[8] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2940_ _0907_ _0598_ _0605_ VGND VGND VPWR VPWR _0606_ sky130_fd_sc_hd__o21a_1
XFILLER_0_29_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2871_ _0529_ _0531_ _1243_ VGND VGND VPWR VPWR _0532_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_29_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_478 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1822_ _0716_ _0796_ _0965_ VGND VGND VPWR VPWR _0966_ sky130_fd_sc_hd__and3_4
X_1753_ _0763_ _0854_ _0897_ VGND VGND VPWR VPWR _0898_ sky130_fd_sc_hd__and3_2
XFILLER_0_13_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1684_ _0828_ _0742_ VGND VGND VPWR VPWR _0829_ sky130_fd_sc_hd__nand2_8
XFILLER_0_20_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2305_ _1003_ _0939_ _0790_ VGND VGND VPWR VPWR _1443_ sky130_fd_sc_hd__and3_2
X_2236_ _1047_ _1374_ _1375_ _0993_ VGND VGND VPWR VPWR _1376_ sky130_fd_sc_hd__a31o_1
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2167_ _1115_ VGND VGND VPWR VPWR _1308_ sky130_fd_sc_hd__buf_4
XFILLER_0_17_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2098_ _1209_ _1218_ _1228_ _1239_ _0843_ _1161_ VGND VGND VPWR VPWR _1240_ sky130_fd_sc_hd__mux4_2
XFILLER_0_48_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3070_ net1 VGND VGND VPWR VPWR _0707_ sky130_fd_sc_hd__buf_4
X_2021_ _1161_ _1162_ VGND VGND VPWR VPWR _1163_ sky130_fd_sc_hd__nor2_1
XFILLER_0_77_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2923_ _0685_ _0585_ _0586_ VGND VGND VPWR VPWR _0587_ sky130_fd_sc_hd__and3_1
XFILLER_0_72_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2854_ _1059_ _0444_ _0944_ VGND VGND VPWR VPWR _0513_ sky130_fd_sc_hd__o21a_1
XFILLER_0_72_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1805_ _0685_ VGND VGND VPWR VPWR _0950_ sky130_fd_sc_hd__buf_4
XFILLER_0_53_470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2785_ _1109_ _0940_ _0928_ _0438_ _1115_ VGND VGND VPWR VPWR _0439_ sky130_fd_sc_hd__o311a_1
X_1736_ _0729_ VGND VGND VPWR VPWR _0881_ sky130_fd_sc_hd__buf_8
XFILLER_0_13_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1667_ _0718_ _0731_ VGND VGND VPWR VPWR _0812_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1598_ _0741_ _0742_ VGND VGND VPWR VPWR _0743_ sky130_fd_sc_hd__nor2_4
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2219_ _0737_ _1041_ _0743_ VGND VGND VPWR VPWR _1359_ sky130_fd_sc_hd__or3_1
XFILLER_0_95_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2570_ _0864_ _1026_ _1065_ VGND VGND VPWR VPWR _0228_ sky130_fd_sc_hd__or3b_1
XFILLER_0_10_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3122_ clknet_2_2__leaf_wb_clk_i _0018_ _0057_ VGND VGND VPWR VPWR weights_inst.data_out\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3053_ net14 _0691_ _0695_ _0699_ VGND VGND VPWR VPWR fsm_inst.next_state\[1\] sky130_fd_sc_hd__o31ai_1
X_2004_ _0835_ _1146_ VGND VGND VPWR VPWR _1147_ sky130_fd_sc_hd__nand2_2
XFILLER_0_77_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2906_ _0956_ _0744_ _1172_ _0568_ _0838_ VGND VGND VPWR VPWR _0569_ sky130_fd_sc_hd__o311a_1
XFILLER_0_60_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2837_ _1322_ _0480_ _0494_ _1242_ VGND VGND VPWR VPWR _0014_ sky130_fd_sc_hd__o211a_1
X_2768_ _0770_ _0340_ _1151_ VGND VGND VPWR VPWR _0422_ sky130_fd_sc_hd__a21o_1
XFILLER_0_41_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1719_ _0833_ VGND VGND VPWR VPWR _0864_ sky130_fd_sc_hd__buf_4
XFILLER_0_41_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2699_ _1180_ _0829_ _1135_ _0963_ VGND VGND VPWR VPWR _0354_ sky130_fd_sc_hd__o31a_1
XTAP_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_495 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_19 _0645_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2622_ _0873_ _0854_ _0739_ VGND VGND VPWR VPWR _0279_ sky130_fd_sc_hd__and3_1
XFILLER_0_23_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2553_ _0936_ _1077_ _0137_ VGND VGND VPWR VPWR _0212_ sky130_fd_sc_hd__or3_1
XFILLER_0_100_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2484_ _1367_ _0886_ _1112_ _1040_ VGND VGND VPWR VPWR _0144_ sky130_fd_sc_hd__a211o_1
X_3105_ clknet_2_3__leaf_wb_clk_i _0023_ _0040_ VGND VGND VPWR VPWR weights_inst.data_out\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3036_ _0684_ VGND VGND VPWR VPWR _0000_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_223 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_340 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput17 wbs_stb_i VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_510 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1984_ _0826_ net54 VGND VGND VPWR VPWR _1127_ sky130_fd_sc_hd__nor2_4
XFILLER_0_70_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2605_ _1342_ _0259_ _0261_ _0843_ VGND VGND VPWR VPWR _0262_ sky130_fd_sc_hd__o211a_1
XFILLER_0_11_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2536_ _0771_ _0983_ VGND VGND VPWR VPWR _0195_ sky130_fd_sc_hd__nor2_1
X_2467_ _1168_ _0076_ _0911_ VGND VGND VPWR VPWR _0128_ sky130_fd_sc_hd__o21a_1
XFILLER_0_47_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2398_ _1003_ _1311_ _1516_ _1109_ VGND VGND VPWR VPWR _0060_ sky130_fd_sc_hd__a211o_1
XFILLER_0_78_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3019_ weights_inst.data_out\[16\] _0666_ VGND VGND VPWR VPWR _0675_ sky130_fd_sc_hd__and2_1
Xwire52 _0773_ VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__buf_4
XFILLER_0_38_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2321_ _0910_ _1175_ _1456_ _1458_ _0685_ VGND VGND VPWR VPWR _1459_ sky130_fd_sc_hd__o311a_1
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2252_ _0729_ _0730_ VGND VGND VPWR VPWR _1391_ sky130_fd_sc_hd__nor2_4
XFILLER_0_85_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2183_ _1188_ _0886_ VGND VGND VPWR VPWR _1323_ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1967_ _0939_ _0797_ VGND VGND VPWR VPWR _1110_ sky130_fd_sc_hd__nand2_2
XFILLER_0_43_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1898_ _1041_ _0996_ _0892_ VGND VGND VPWR VPWR _1042_ sky130_fd_sc_hd__and3_2
XFILLER_0_31_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2519_ _1158_ _0151_ _0178_ _1242_ VGND VGND VPWR VPWR _0006_ sky130_fd_sc_hd__o211a_1
XFILLER_0_59_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold6 net10 VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2870_ _1403_ _1379_ _0124_ _0530_ _1308_ VGND VGND VPWR VPWR _0531_ sky130_fd_sc_hd__o311a_1
XFILLER_0_29_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1821_ _0729_ _0731_ _0795_ VGND VGND VPWR VPWR _0965_ sky130_fd_sc_hd__a21o_4
XFILLER_0_13_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1752_ _0742_ _0896_ VGND VGND VPWR VPWR _0897_ sky130_fd_sc_hd__nand2_1
X_1683_ _0795_ VGND VGND VPWR VPWR _0828_ sky130_fd_sc_hd__buf_8
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_73 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2304_ _0993_ _1431_ _1435_ _1437_ _1441_ VGND VGND VPWR VPWR _1442_ sky130_fd_sc_hd__o32a_1
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2235_ _1124_ _1221_ _1097_ _0878_ _0922_ VGND VGND VPWR VPWR _1375_ sky130_fd_sc_hd__a221o_1
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2166_ _1306_ _1056_ _1107_ VGND VGND VPWR VPWR _1307_ sky130_fd_sc_hd__or3b_4
X_2097_ _1198_ _1231_ _1234_ _1238_ VGND VGND VPWR VPWR _1239_ sky130_fd_sc_hd__a31o_1
XFILLER_0_63_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2999_ _0662_ VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__buf_1
XFILLER_0_28_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2020_ _0825_ _0918_ _0802_ VGND VGND VPWR VPWR _1162_ sky130_fd_sc_hd__and3_2
XFILLER_0_89_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2922_ _1265_ _1334_ _0984_ VGND VGND VPWR VPWR _0586_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_85_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2853_ _0734_ _1146_ _1167_ _0511_ _1178_ VGND VGND VPWR VPWR _0512_ sky130_fd_sc_hd__a311o_1
XFILLER_0_45_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2784_ _1491_ _1016_ _1022_ _1211_ VGND VGND VPWR VPWR _0438_ sky130_fd_sc_hd__o31ai_1
X_1804_ _0947_ _0948_ VGND VGND VPWR VPWR _0949_ sky130_fd_sc_hd__nand2_1
X_1735_ _0828_ _0711_ VGND VGND VPWR VPWR _0880_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_53_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1666_ _0810_ VGND VGND VPWR VPWR _0811_ sky130_fd_sc_hd__buf_4
X_1597_ _0711_ VGND VGND VPWR VPWR _0742_ sky130_fd_sc_hd__buf_8
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2218_ _1123_ _0797_ _0785_ VGND VGND VPWR VPWR _1358_ sky130_fd_sc_hd__a21o_1
XFILLER_0_95_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2149_ _0725_ _1288_ _1289_ _1022_ _1187_ VGND VGND VPWR VPWR _1290_ sky130_fd_sc_hd__o32a_1
XFILLER_0_95_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_438 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_279 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3121_ clknet_2_3__leaf_wb_clk_i _0017_ _0056_ VGND VGND VPWR VPWR weights_inst.data_out\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3052_ fsm_inst.current_state\[1\] fsm_inst.current_state\[0\] VGND VGND VPWR VPWR
+ _0699_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2003_ _0828_ _0758_ VGND VGND VPWR VPWR _1146_ sky130_fd_sc_hd__nand2_2
XFILLER_0_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2905_ _0802_ _1105_ _1324_ _0892_ _0834_ VGND VGND VPWR VPWR _0568_ sky130_fd_sc_hd__a221o_1
XFILLER_0_45_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2836_ _1365_ _0492_ _0493_ _1322_ VGND VGND VPWR VPWR _0494_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_5_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2767_ _0817_ _1077_ _1410_ _1050_ _0985_ VGND VGND VPWR VPWR _0421_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_77_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1718_ net70 VGND VGND VPWR VPWR _0863_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_41_474 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2698_ _0755_ _1167_ VGND VGND VPWR VPWR _0353_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_187 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1649_ _0742_ _0793_ VGND VGND VPWR VPWR _0794_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_327 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2621_ _1199_ _1506_ _0080_ VGND VGND VPWR VPWR _0278_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_2_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2552_ _1403_ _1300_ _0209_ _0210_ _1356_ VGND VGND VPWR VPWR _0211_ sky130_fd_sc_hd__o311a_1
XFILLER_0_23_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_271 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2483_ _1356_ _0139_ _0142_ VGND VGND VPWR VPWR _0143_ sky130_fd_sc_hd__o21ba_1
X_3104_ clknet_2_0__leaf_wb_clk_i _0022_ _0039_ VGND VGND VPWR VPWR weights_inst.data_out\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_3035_ fsm_inst.current_state\[1\] fsm_inst.current_state\[0\] fsm_inst.current_state\[2\]
+ VGND VGND VPWR VPWR _0684_ sky130_fd_sc_hd__and3b_1
XFILLER_0_77_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2819_ _0878_ _1213_ _0450_ _1140_ VGND VGND VPWR VPWR _0476_ sky130_fd_sc_hd__a211o_1
XFILLER_0_14_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput18 wbs_we_i VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__buf_1
XFILLER_0_52_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1983_ _1124_ _1106_ _1125_ _1060_ VGND VGND VPWR VPWR _1126_ sky130_fd_sc_hd__a211o_1
XFILLER_0_43_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2604_ _1256_ _1214_ _0257_ _0260_ _0915_ VGND VGND VPWR VPWR _0261_ sky130_fd_sc_hd__a311o_1
XFILLER_0_11_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2535_ _0861_ _0185_ _0192_ _0193_ VGND VGND VPWR VPWR _0194_ sky130_fd_sc_hd__o31a_1
X_2466_ _1273_ _0123_ _0126_ VGND VGND VPWR VPWR _0127_ sky130_fd_sc_hd__or3_1
X_2397_ _1532_ _1350_ _0752_ VGND VGND VPWR VPWR _0059_ sky130_fd_sc_hd__a21o_1
XFILLER_0_78_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3018_ _0674_ VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__buf_1
XFILLER_0_78_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2320_ _0723_ _1066_ _1457_ VGND VGND VPWR VPWR _1458_ sky130_fd_sc_hd__or3_1
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2251_ _0892_ _0973_ _1324_ _1267_ _1040_ VGND VGND VPWR VPWR _1390_ sky130_fd_sc_hd__a311o_1
X_2182_ _0863_ VGND VGND VPWR VPWR _1322_ sky130_fd_sc_hd__buf_2
XFILLER_0_75_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1966_ _0944_ VGND VGND VPWR VPWR _1109_ sky130_fd_sc_hd__buf_4
XFILLER_0_7_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1897_ _0826_ VGND VGND VPWR VPWR _1041_ sky130_fd_sc_hd__buf_4
XFILLER_0_101_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2518_ _1197_ _0177_ VGND VGND VPWR VPWR _0178_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2449_ _1117_ _0813_ _0867_ VGND VGND VPWR VPWR _0110_ sky130_fd_sc_hd__or3_1
XFILLER_0_75_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold7 _0858_ VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_89_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1820_ _0834_ VGND VGND VPWR VPWR _0964_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_13_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1751_ _0717_ _0708_ VGND VGND VPWR VPWR _0896_ sky130_fd_sc_hd__nor2_8
XFILLER_0_52_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1682_ _0825_ _0826_ _0746_ VGND VGND VPWR VPWR _0827_ sky130_fd_sc_hd__and3_4
XFILLER_0_21_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2303_ _0963_ _1440_ _0993_ VGND VGND VPWR VPWR _1441_ sky130_fd_sc_hd__o21ai_1
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2234_ _1229_ _0965_ _1059_ net56 _1140_ VGND VGND VPWR VPWR _1374_ sky130_fd_sc_hd__a221o_1
X_2165_ _0891_ _0972_ _0768_ VGND VGND VPWR VPWR _1306_ sky130_fd_sc_hd__a21oi_1
X_2096_ _1235_ _0912_ _0980_ _1237_ _0950_ VGND VGND VPWR VPWR _1238_ sky130_fd_sc_hd__o311a_1
XFILLER_0_48_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2998_ weights_inst.data_out\[6\] _0654_ VGND VGND VPWR VPWR _0662_ sky130_fd_sc_hd__and2_1
XFILLER_0_71_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1949_ _1089_ _0769_ _0713_ _1091_ VGND VGND VPWR VPWR _1092_ sky130_fd_sc_hd__a31o_1
XFILLER_0_16_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2921_ _0833_ _0768_ _0965_ VGND VGND VPWR VPWR _0585_ sky130_fd_sc_hd__or3_1
XFILLER_0_57_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2852_ _0827_ _0105_ _1180_ VGND VGND VPWR VPWR _0511_ sky130_fd_sc_hd__o21a_1
X_1803_ _0926_ _0930_ VGND VGND VPWR VPWR _0948_ sky130_fd_sc_hd__nor2_8
X_2783_ _0426_ _0436_ _0849_ VGND VGND VPWR VPWR _0437_ sky130_fd_sc_hd__o21ai_4
X_1734_ _0878_ _0813_ VGND VGND VPWR VPWR _0879_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1665_ _0799_ VGND VGND VPWR VPWR _0810_ sky130_fd_sc_hd__buf_4
XFILLER_0_21_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1596_ _0708_ VGND VGND VPWR VPWR _0741_ sky130_fd_sc_hd__clkbuf_8
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2217_ _0752_ _1190_ _1354_ _1355_ _1356_ VGND VGND VPWR VPWR _1357_ sky130_fd_sc_hd__o311ai_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2148_ _1123_ _0971_ _1136_ VGND VGND VPWR VPWR _1289_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_95_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2079_ _0757_ _0804_ VGND VGND VPWR VPWR _1221_ sky130_fd_sc_hd__nor2_4
XFILLER_0_76_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3120_ clknet_2_2__leaf_wb_clk_i _0016_ _0055_ VGND VGND VPWR VPWR weights_inst.data_out\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3051_ _0688_ _0691_ _0695_ _0698_ VGND VGND VPWR VPWR fsm_inst.next_state\[0\] sky130_fd_sc_hd__o31ai_1
XFILLER_0_26_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2002_ _1140_ _1141_ _1142_ _1144_ VGND VGND VPWR VPWR _1145_ sky130_fd_sc_hd__o31a_1
XFILLER_0_77_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2904_ _0824_ _1106_ _0358_ VGND VGND VPWR VPWR _0567_ sky130_fd_sc_hd__a21o_1
X_2835_ _0917_ _1379_ _0270_ _1161_ VGND VGND VPWR VPWR _0493_ sky130_fd_sc_hd__a211o_1
XFILLER_0_14_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2766_ _1299_ _0076_ _0418_ _0801_ _1115_ VGND VGND VPWR VPWR _0419_ sky130_fd_sc_hd__o221a_1
XFILLER_0_13_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1717_ _0845_ _0846_ _0847_ VGND VGND VPWR VPWR _0862_ sky130_fd_sc_hd__and3_1
XFILLER_0_5_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2697_ _1347_ _1254_ net51 _0655_ VGND VGND VPWR VPWR _0352_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_41_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1648_ _0717_ _0708_ VGND VGND VPWR VPWR _0793_ sky130_fd_sc_hd__or2b_1
XFILLER_0_1_594 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1579_ _0723_ VGND VGND VPWR VPWR _0724_ sky130_fd_sc_hd__buf_4
XTAP_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_339 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2620_ _1250_ _0272_ _0276_ VGND VGND VPWR VPWR _0277_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_88_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2551_ _1367_ _0886_ _0961_ _0829_ _1264_ VGND VGND VPWR VPWR _0210_ sky130_fd_sc_hd__a221o_1
XFILLER_0_10_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_283 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2482_ _0957_ _0767_ _0890_ _0141_ _0778_ VGND VGND VPWR VPWR _0142_ sky130_fd_sc_hd__o311a_1
X_3103_ clknet_2_0__leaf_wb_clk_i _0021_ _0038_ VGND VGND VPWR VPWR weights_inst.data_out\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_3034_ _0683_ VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__buf_2
XFILLER_0_37_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2818_ _0472_ _0474_ VGND VGND VPWR VPWR _0475_ sky130_fd_sc_hd__xnor2_1
X_2749_ _0917_ _1045_ _1189_ _0957_ VGND VGND VPWR VPWR _0403_ sky130_fd_sc_hd__a211o_1
XFILLER_0_41_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1982_ _0769_ _0802_ VGND VGND VPWR VPWR _1125_ sky130_fd_sc_hd__nor2_2
XFILLER_0_7_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2603_ _0869_ _1236_ _1399_ _0770_ _0810_ VGND VGND VPWR VPWR _0260_ sky130_fd_sc_hd__o221a_1
XFILLER_0_30_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2534_ _0645_ _1050_ _0146_ VGND VGND VPWR VPWR _0193_ sky130_fd_sc_hd__or3_1
XFILLER_0_11_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2465_ _1335_ _0124_ _1457_ _0125_ _1278_ VGND VGND VPWR VPWR _0126_ sky130_fd_sc_hd__o311a_1
X_2396_ _0947_ _0931_ VGND VGND VPWR VPWR _1532_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3017_ weights_inst.data_out\[15\] _0666_ VGND VGND VPWR VPWR _0674_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2250_ _0786_ _1031_ _0875_ VGND VGND VPWR VPWR _1389_ sky130_fd_sc_hd__a21o_1
X_2181_ _1158_ _1163_ _1272_ _1321_ _0859_ VGND VGND VPWR VPWR _0022_ sky130_fd_sc_hd__o311a_1
X_1965_ _0645_ _1102_ _1104_ _1107_ _0848_ VGND VGND VPWR VPWR _1108_ sky130_fd_sc_hd__a221o_1
XFILLER_0_50_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1896_ _1028_ VGND VGND VPWR VPWR _1040_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_70_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2517_ _0157_ _0162_ _0169_ _0176_ _0843_ _0645_ VGND VGND VPWR VPWR _0177_ sky130_fd_sc_hd__mux4_2
X_2448_ _1120_ net56 VGND VGND VPWR VPWR _0109_ sky130_fd_sc_hd__nor2_1
XFILLER_0_52_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2379_ _0975_ _0924_ _0851_ VGND VGND VPWR VPWR _1516_ sky130_fd_sc_hd__and3_1
XFILLER_0_75_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold8 _1157_ VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1750_ _0889_ _0890_ _0894_ VGND VGND VPWR VPWR _0895_ sky130_fd_sc_hd__o21a_1
XFILLER_0_20_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1681_ _0763_ VGND VGND VPWR VPWR _0826_ sky130_fd_sc_hd__buf_4
XFILLER_0_96_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2302_ _0964_ _1438_ _1439_ _1292_ _0900_ VGND VGND VPWR VPWR _1440_ sky130_fd_sc_hd__o32a_1
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2233_ _1180_ _0988_ _1200_ VGND VGND VPWR VPWR _1373_ sky130_fd_sc_hd__or3_1
X_2164_ _0826_ _0989_ VGND VGND VPWR VPWR _1305_ sky130_fd_sc_hd__nor2_2
XFILLER_0_45_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2095_ _0929_ _0960_ _1236_ _0956_ VGND VGND VPWR VPWR _1237_ sky130_fd_sc_hd__a211o_1
XFILLER_0_75_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2997_ _0660_ VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__buf_1
X_1948_ _0723_ _1090_ VGND VGND VPWR VPWR _1091_ sky130_fd_sc_hd__or2_1
XFILLER_0_71_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1879_ _0820_ net52 VGND VGND VPWR VPWR _1023_ sky130_fd_sc_hd__nor2_4
XFILLER_0_9_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_451 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2920_ _0799_ _1466_ _0075_ _0583_ _0776_ VGND VGND VPWR VPWR _0584_ sky130_fd_sc_hd__o311a_1
XFILLER_0_57_245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2851_ _1250_ _0508_ _0509_ VGND VGND VPWR VPWR _0510_ sky130_fd_sc_hd__nand3_1
XFILLER_0_57_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2782_ _0952_ _0428_ _0430_ _0435_ _0645_ VGND VGND VPWR VPWR _0436_ sky130_fd_sc_hd__o311a_1
X_1802_ _0897_ VGND VGND VPWR VPWR _0947_ sky130_fd_sc_hd__buf_4
X_1733_ _0877_ VGND VGND VPWR VPWR _0878_ sky130_fd_sc_hd__buf_6
XFILLER_0_5_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1664_ _0798_ _0801_ _0808_ VGND VGND VPWR VPWR _0809_ sky130_fd_sc_hd__or3b_1
XFILLER_0_0_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1595_ _0727_ VGND VGND VPWR VPWR _0740_ sky130_fd_sc_hd__clkbuf_8
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2216_ _0782_ VGND VGND VPWR VPWR _1356_ sky130_fd_sc_hd__clkbuf_4
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2147_ _1117_ _0854_ _0927_ VGND VGND VPWR VPWR _1288_ sky130_fd_sc_hd__and3_2
XFILLER_0_95_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2078_ _0944_ _1016_ VGND VGND VPWR VPWR _1220_ sky130_fd_sc_hd__nor2_1
XFILLER_0_72_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3050_ fsm_inst.current_state\[0\] _0697_ _0693_ VGND VGND VPWR VPWR _0698_ sky130_fd_sc_hd__a21bo_1
X_2001_ _0798_ _1143_ _1060_ VGND VGND VPWR VPWR _1144_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_89_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2903_ _0721_ _0739_ _1072_ _1159_ _0956_ VGND VGND VPWR VPWR _0566_ sky130_fd_sc_hd__a221o_1
XFILLER_0_58_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2834_ _1164_ _0482_ _0485_ _0488_ _0491_ VGND VGND VPWR VPWR _0492_ sky130_fd_sc_hd__o32a_1
XFILLER_0_14_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2765_ _0805_ _0417_ _1095_ VGND VGND VPWR VPWR _0418_ sky130_fd_sc_hd__o21a_1
XFILLER_0_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1716_ _0860_ VGND VGND VPWR VPWR _0861_ sky130_fd_sc_hd__clkbuf_4
X_2696_ _1243_ _0343_ _0350_ _0655_ VGND VGND VPWR VPWR _0351_ sky130_fd_sc_hd__o211a_1
XFILLER_0_1_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1647_ _0789_ _0791_ VGND VGND VPWR VPWR _0792_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1578_ _0473_ _0505_ VGND VGND VPWR VPWR _0723_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_6_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2550_ _0758_ _0976_ VGND VGND VPWR VPWR _0209_ sky130_fd_sc_hd__and2_2
XFILLER_0_50_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2481_ _1245_ _0140_ _0873_ VGND VGND VPWR VPWR _0141_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_50_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3102_ clknet_2_0__leaf_wb_clk_i _0019_ _0037_ VGND VGND VPWR VPWR weights_inst.data_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_3033_ weights_inst.data_out\[23\] net55 VGND VGND VPWR VPWR _0683_ sky130_fd_sc_hd__and2_1
XFILLER_0_77_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2817_ _0936_ _1399_ VGND VGND VPWR VPWR _0474_ sky130_fd_sc_hd__nand2_1
X_2748_ _0929_ _1206_ VGND VGND VPWR VPWR _0402_ sky130_fd_sc_hd__nand2_1
X_2679_ _1298_ _0326_ _0328_ _0334_ _1039_ VGND VGND VPWR VPWR _0335_ sky130_fd_sc_hd__o311a_1
XFILLER_0_96_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1981_ _1123_ VGND VGND VPWR VPWR _1124_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_99_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2602_ _0811_ _1160_ _0256_ _0257_ _0258_ VGND VGND VPWR VPWR _0259_ sky130_fd_sc_hd__a32o_1
X_2533_ _0187_ _0188_ _0191_ VGND VGND VPWR VPWR _0192_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_23_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2464_ _1063_ _1053_ _1277_ VGND VGND VPWR VPWR _0125_ sky130_fd_sc_hd__or3_1
X_2395_ _1256_ _1233_ _1530_ VGND VGND VPWR VPWR _1531_ sky130_fd_sc_hd__or3_1
XFILLER_0_48_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3016_ _0672_ VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__buf_1
XFILLER_0_93_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire55 net88 VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_93_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2180_ _1297_ _1320_ _1197_ VGND VGND VPWR VPWR _1321_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_75_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1964_ _0817_ _1106_ VGND VGND VPWR VPWR _1107_ sky130_fd_sc_hd__nand2_2
XFILLER_0_70_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1895_ _0860_ VGND VGND VPWR VPWR _1039_ sky130_fd_sc_hd__buf_4
XFILLER_0_70_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2516_ _1198_ _0170_ _0171_ _0175_ VGND VGND VPWR VPWR _0176_ sky130_fd_sc_hd__a31o_1
X_2447_ _1250_ _0103_ _0104_ _0107_ _1273_ VGND VGND VPWR VPWR _0108_ sky130_fd_sc_hd__a311o_1
XFILLER_0_45_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2378_ _1012_ _1347_ _1202_ _1291_ VGND VGND VPWR VPWR _1515_ sky130_fd_sc_hd__a211o_1
XFILLER_0_78_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold9 wbs_adr_i[7] VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1680_ _0793_ VGND VGND VPWR VPWR _0825_ sky130_fd_sc_hd__buf_6
XFILLER_0_21_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2301_ _0716_ _0829_ net56 VGND VGND VPWR VPWR _1439_ sky130_fd_sc_hd__and3_1
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2232_ _0917_ _1066_ _0940_ _1165_ VGND VGND VPWR VPWR _1372_ sky130_fd_sc_hd__a211o_1
X_2163_ _1299_ _1300_ _1302_ _1303_ _0779_ VGND VGND VPWR VPWR _1304_ sky130_fd_sc_hd__o311a_1
X_2094_ _0828_ _0866_ VGND VGND VPWR VPWR _1236_ sky130_fd_sc_hd__nor2_4
XFILLER_0_45_75 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2996_ weights_inst.data_out\[5\] _0654_ VGND VGND VPWR VPWR _0660_ sky130_fd_sc_hd__and2_1
XFILLER_0_71_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1947_ _0763_ _0999_ VGND VGND VPWR VPWR _1090_ sky130_fd_sc_hd__nor2_1
XFILLER_0_71_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1878_ _1012_ _0970_ VGND VGND VPWR VPWR _1022_ sky130_fd_sc_hd__nor2_2
XFILLER_0_31_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2850_ _0917_ _0807_ _1389_ VGND VGND VPWR VPWR _0509_ sky130_fd_sc_hd__a21o_1
XFILLER_0_57_257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1801_ _0708_ _0710_ VGND VGND VPWR VPWR _0946_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_38_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2781_ _1047_ _0431_ _0432_ _0434_ _0993_ VGND VGND VPWR VPWR _0435_ sky130_fd_sc_hd__a311o_1
X_1732_ _0757_ VGND VGND VPWR VPWR _0877_ sky130_fd_sc_hd__buf_6
X_1663_ _0803_ _0807_ VGND VGND VPWR VPWR _0808_ sky130_fd_sc_hd__nand2_1
X_1594_ _0738_ VGND VGND VPWR VPWR _0739_ sky130_fd_sc_hd__clkbuf_8
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2215_ _0971_ _1079_ _1330_ _0911_ VGND VGND VPWR VPWR _1355_ sky130_fd_sc_hd__a211o_1
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2146_ _0963_ VGND VGND VPWR VPWR _1287_ sky130_fd_sc_hd__clkbuf_4
X_2077_ _0924_ VGND VGND VPWR VPWR _1219_ sky130_fd_sc_hd__buf_4
XFILLER_0_76_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2979_ _1356_ _0646_ _0647_ _0617_ VGND VGND VPWR VPWR _0648_ sky130_fd_sc_hd__a31o_1
XFILLER_0_44_441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2000_ _1003_ _0926_ _0823_ VGND VGND VPWR VPWR _1143_ sky130_fd_sc_hd__and3_1
XFILLER_0_58_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2902_ _0934_ _0562_ _0563_ _0564_ VGND VGND VPWR VPWR _0565_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_85_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2833_ _1356_ _0489_ _0490_ _0952_ VGND VGND VPWR VPWR _0491_ sky130_fd_sc_hd__a31o_1
XFILLER_0_5_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2764_ _0975_ _1113_ VGND VGND VPWR VPWR _0417_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1715_ _0602_ _0623_ VGND VGND VPWR VPWR _0860_ sky130_fd_sc_hd__xor2_4
X_2695_ _0347_ _0349_ _1243_ VGND VGND VPWR VPWR _0350_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_1_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1646_ _0727_ _0790_ VGND VGND VPWR VPWR _0791_ sky130_fd_sc_hd__nand2_4
X_1577_ _0713_ _0721_ VGND VGND VPWR VPWR _0722_ sky130_fd_sc_hd__nand2_4
XFILLER_0_67_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2129_ _0783_ _1260_ _1263_ _1269_ VGND VGND VPWR VPWR _1270_ sky130_fd_sc_hd__a31o_1
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2480_ _0787_ _0813_ VGND VGND VPWR VPWR _0140_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3101_ clknet_2_1__leaf_wb_clk_i _0015_ _0036_ VGND VGND VPWR VPWR weights_inst.data_out\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_3032_ _0682_ VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__buf_1
XFILLER_0_77_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2816_ _0916_ _1077_ _1023_ VGND VGND VPWR VPWR _0472_ sky130_fd_sc_hd__a21o_1
XFILLER_0_14_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2747_ _0655_ _0400_ VGND VGND VPWR VPWR _0401_ sky130_fd_sc_hd__nor2_1
XFILLER_0_75_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2678_ _1287_ _0329_ _0330_ _0333_ _1318_ VGND VGND VPWR VPWR _0334_ sky130_fd_sc_hd__a311o_1
XFILLER_0_78_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1629_ _0770_ net52 VGND VGND VPWR VPWR _0774_ sky130_fd_sc_hd__nor2_2
XFILLER_0_1_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1980_ _0741_ VGND VGND VPWR VPWR _1123_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_67_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_311 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2601_ _0751_ _0928_ VGND VGND VPWR VPWR _0258_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2532_ _0703_ _0189_ _0190_ _1193_ VGND VGND VPWR VPWR _0191_ sky130_fd_sc_hd__a31o_1
XFILLER_0_51_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2463_ _1011_ _0903_ VGND VGND VPWR VPWR _0124_ sky130_fd_sc_hd__nor2_4
X_2394_ _0785_ _0713_ _0959_ VGND VGND VPWR VPWR _1530_ sky130_fd_sc_hd__and3_1
XFILLER_0_48_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3015_ weights_inst.data_out\[14\] _0666_ VGND VGND VPWR VPWR _0672_ sky130_fd_sc_hd__and2_1
XFILLER_0_64_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1963_ _1105_ VGND VGND VPWR VPWR _1106_ sky130_fd_sc_hd__buf_4
X_1894_ _0995_ _1037_ _0849_ VGND VGND VPWR VPWR _1038_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_55_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2515_ _1235_ _1127_ _1162_ _0174_ _0950_ VGND VGND VPWR VPWR _0175_ sky130_fd_sc_hd__o311a_1
X_2446_ _1291_ net51 _1443_ _0106_ _0703_ VGND VGND VPWR VPWR _0107_ sky130_fd_sc_hd__o311a_1
XFILLER_0_75_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2377_ _1281_ _1491_ _1511_ _1513_ _1310_ VGND VGND VPWR VPWR _1514_ sky130_fd_sc_hd__o311a_1
XFILLER_0_78_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2300_ _0877_ _0903_ VGND VGND VPWR VPWR _1438_ sky130_fd_sc_hd__nor2_1
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2231_ _0752_ _1182_ _1277_ _1370_ _1356_ VGND VGND VPWR VPWR _1371_ sky130_fd_sc_hd__o311a_1
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2162_ _1000_ _1043_ _1020_ _1301_ _1180_ VGND VGND VPWR VPWR _1303_ sky130_fd_sc_hd__a221o_1
XFILLER_0_45_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2093_ _0835_ VGND VGND VPWR VPWR _1235_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_88_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2995_ _0659_ VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__buf_1
XFILLER_0_44_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1946_ _0772_ VGND VGND VPWR VPWR _1089_ sky130_fd_sc_hd__buf_4
XFILLER_0_28_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1877_ _0786_ _1019_ _0807_ _1020_ _0755_ VGND VGND VPWR VPWR _1021_ sky130_fd_sc_hd__a221o_1
XFILLER_0_16_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2429_ _0999_ _1221_ _1112_ _1219_ _0910_ VGND VGND VPWR VPWR _0091_ sky130_fd_sc_hd__a221o_1
XFILLER_0_79_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1800_ _0944_ VGND VGND VPWR VPWR _0945_ sky130_fd_sc_hd__buf_4
XFILLER_0_26_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2780_ _1225_ _1330_ _0433_ _0777_ VGND VGND VPWR VPWR _0434_ sky130_fd_sc_hd__o211a_2
XFILLER_0_53_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1731_ _0815_ _0817_ VGND VGND VPWR VPWR _0876_ sky130_fd_sc_hd__nand2_1
X_1662_ _0806_ VGND VGND VPWR VPWR _0807_ sky130_fd_sc_hd__buf_4
XFILLER_0_21_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1593_ _0735_ _0737_ VGND VGND VPWR VPWR _0738_ sky130_fd_sc_hd__nand2_4
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2214_ _0926_ _0790_ _0947_ VGND VGND VPWR VPWR _1354_ sky130_fd_sc_hd__and3_4
X_2145_ _1281_ _1265_ _1282_ _1284_ _1285_ VGND VGND VPWR VPWR _1286_ sky130_fd_sc_hd__o311a_1
XFILLER_0_76_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2076_ _1178_ _1210_ _1212_ _1217_ VGND VGND VPWR VPWR _1218_ sky130_fd_sc_hd__a31o_1
XFILLER_0_76_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2978_ _0983_ _0931_ _1300_ _0923_ VGND VGND VPWR VPWR _0647_ sky130_fd_sc_hd__a211o_1
XFILLER_0_71_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1929_ _0765_ net74 VGND VGND VPWR VPWR _1073_ sky130_fd_sc_hd__nand2_8
XFILLER_0_44_453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_103 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2901_ _0561_ _1329_ VGND VGND VPWR VPWR _0564_ sky130_fd_sc_hd__or2b_1
XFILLER_0_58_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2832_ _1232_ _1367_ _0867_ _1152_ _0801_ VGND VGND VPWR VPWR _0490_ sky130_fd_sc_hd__a311o_1
X_2763_ _0734_ _0856_ _0415_ _0703_ VGND VGND VPWR VPWR _0416_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_5_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1714_ net66 VGND VGND VPWR VPWR _0859_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_53_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2694_ _1403_ _0948_ _1002_ _0348_ _1308_ VGND VGND VPWR VPWR _0349_ sky130_fd_sc_hd__o311a_1
X_1645_ _0708_ _0731_ VGND VGND VPWR VPWR _0790_ sky130_fd_sc_hd__nand2_4
X_1576_ _0716_ _0720_ VGND VGND VPWR VPWR _0721_ sky130_fd_sc_hd__nor2_4
XFILLER_0_21_191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2128_ _1264_ _1265_ _1266_ _1268_ _1047_ VGND VGND VPWR VPWR _1269_ sky130_fd_sc_hd__o311a_1
X_2059_ _1199_ _1014_ _1200_ _1056_ VGND VGND VPWR VPWR _1201_ sky130_fd_sc_hd__a211o_1
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3100_ clknet_2_0__leaf_wb_clk_i _0004_ _0035_ VGND VGND VPWR VPWR weights_inst.data_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3031_ weights_inst.data_out\[22\] net55 VGND VGND VPWR VPWR _0682_ sky130_fd_sc_hd__and2_1
XFILLER_0_37_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2815_ _1281_ _0990_ _1470_ _0470_ _1308_ VGND VGND VPWR VPWR _0471_ sky130_fd_sc_hd__o311a_1
XFILLER_0_61_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2746_ _0673_ _0392_ _0394_ _0396_ _0399_ VGND VGND VPWR VPWR _0400_ sky130_fd_sc_hd__o32a_1
XFILLER_0_14_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2677_ _0945_ _0747_ _1027_ _0332_ _0778_ VGND VGND VPWR VPWR _0333_ sky130_fd_sc_hd__o311a_1
XFILLER_0_68_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1628_ _0729_ _0771_ _0772_ VGND VGND VPWR VPWR _0773_ sky130_fd_sc_hd__a21oi_1
X_1559_ _0473_ _0495_ _0484_ VGND VGND VPWR VPWR _0679_ sky130_fd_sc_hd__a21boi_4
XFILLER_0_94_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2600_ _0715_ _0998_ _0818_ VGND VGND VPWR VPWR _0257_ sky130_fd_sc_hd__or3_2
XFILLER_0_23_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2531_ _1083_ _0827_ _0154_ VGND VGND VPWR VPWR _0190_ sky130_fd_sc_hd__or3_1
XFILLER_0_51_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2462_ _1291_ _1448_ _1511_ _0122_ _1198_ VGND VGND VPWR VPWR _0123_ sky130_fd_sc_hd__o311a_1
X_2393_ _1158_ _1496_ _1529_ _1242_ VGND VGND VPWR VPWR _0026_ sky130_fd_sc_hd__o211a_1
XFILLER_0_64_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3014_ _0671_ VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__buf_1
XFILLER_0_64_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2729_ _1252_ _1334_ _0752_ VGND VGND VPWR VPWR _0383_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_100_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1962_ _0727_ _0813_ VGND VGND VPWR VPWR _1105_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1893_ _1006_ _1018_ _1035_ _1036_ VGND VGND VPWR VPWR _1037_ sky130_fd_sc_hd__o211a_1
XFILLER_0_43_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2514_ _1136_ _0172_ _0173_ _0956_ VGND VGND VPWR VPWR _0174_ sky130_fd_sc_hd__a211o_1
XFILLER_0_59_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2445_ _1049_ _1079_ _0105_ VGND VGND VPWR VPWR _0106_ sky130_fd_sc_hd__or3_1
X_2376_ _1512_ _0725_ _0761_ VGND VGND VPWR VPWR _1513_ sky130_fd_sc_hd__or3b_1
XFILLER_0_91_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2230_ _0945_ _0733_ _1305_ VGND VGND VPWR VPWR _1370_ sky130_fd_sc_hd__or3_1
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2161_ _1089_ _1301_ VGND VGND VPWR VPWR _1302_ sky130_fd_sc_hd__and2_2
X_2092_ _0942_ _1233_ VGND VGND VPWR VPWR _1234_ sky130_fd_sc_hd__or2_1
XFILLER_0_88_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2994_ weights_inst.data_out\[4\] _0654_ VGND VGND VPWR VPWR _0659_ sky130_fd_sc_hd__and2_1
X_1945_ _0771_ _0825_ VGND VGND VPWR VPWR _1088_ sky130_fd_sc_hd__nor2_4
XFILLER_0_44_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1876_ _0831_ VGND VGND VPWR VPWR _1020_ sky130_fd_sc_hd__buf_4
XFILLER_0_3_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2428_ _0088_ _0089_ _1278_ VGND VGND VPWR VPWR _0090_ sky130_fd_sc_hd__a21oi_1
X_2359_ _1365_ _1481_ _1495_ VGND VGND VPWR VPWR _1496_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_98_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_418 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1730_ _0754_ VGND VGND VPWR VPWR _0875_ sky130_fd_sc_hd__buf_4
X_1661_ _0740_ _0805_ VGND VGND VPWR VPWR _0806_ sky130_fd_sc_hd__nor2_8
XFILLER_0_40_159 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1592_ _0736_ VGND VGND VPWR VPWR _0737_ sky130_fd_sc_hd__buf_8
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2213_ _1342_ _1346_ _1349_ _1352_ _0673_ VGND VGND VPWR VPWR _1353_ sky130_fd_sc_hd__o311a_1
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2144_ _0978_ VGND VGND VPWR VPWR _1285_ sky130_fd_sc_hd__buf_4
XFILLER_0_56_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2075_ _1063_ _1099_ _1152_ _1216_ _0950_ VGND VGND VPWR VPWR _1217_ sky130_fd_sc_hd__o311a_1
XFILLER_0_76_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2977_ _1347_ _0787_ _1206_ _0911_ VGND VGND VPWR VPWR _0646_ sky130_fd_sc_hd__a211o_1
XFILLER_0_44_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1928_ _0784_ _1031_ VGND VGND VPWR VPWR _1072_ sky130_fd_sc_hd__nor2_8
XFILLER_0_44_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1859_ _0794_ VGND VGND VPWR VPWR _1003_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_31_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_476 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2900_ _0944_ _0948_ _1433_ _0777_ VGND VGND VPWR VPWR _0563_ sky130_fd_sc_hd__o31a_1
XFILLER_0_58_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2831_ _1343_ _1019_ _0971_ _1189_ _0911_ VGND VGND VPWR VPWR _0489_ sky130_fd_sc_hd__a311o_1
XFILLER_0_26_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2762_ _1219_ _1023_ _0762_ VGND VGND VPWR VPWR _0415_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_26_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1713_ net8 net9 net65 VGND VGND VPWR VPWR _0858_ sky130_fd_sc_hd__o21ai_1
X_2693_ _1000_ _0816_ _1023_ _1219_ _1264_ VGND VGND VPWR VPWR _0348_ sky130_fd_sc_hd__a221o_1
XFILLER_0_13_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1644_ _0786_ _0788_ _0755_ VGND VGND VPWR VPWR _0789_ sky130_fd_sc_hd__o21a_1
X_1575_ _0711_ _0719_ VGND VGND VPWR VPWR _0720_ sky130_fd_sc_hd__nor2_4
XTAP_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2127_ _1011_ _0739_ _0937_ _1267_ _1083_ VGND VGND VPWR VPWR _1268_ sky130_fd_sc_hd__a311o_1
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2058_ _0852_ _1015_ _0851_ VGND VGND VPWR VPWR _1200_ sky130_fd_sc_hd__and3_4
XFILLER_0_76_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_476 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3030_ _0681_ VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__buf_1
XFILLER_0_53_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2814_ _1347_ _0973_ _0214_ _0923_ VGND VGND VPWR VPWR _0470_ sky130_fd_sc_hd__a211o_1
X_2745_ _1342_ _0397_ _0398_ _0952_ VGND VGND VPWR VPWR _0399_ sky130_fd_sc_hd__a31o_1
XFILLER_0_78_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2676_ _1136_ _0854_ _1325_ _0331_ _0750_ VGND VGND VPWR VPWR _0332_ sky130_fd_sc_hd__a311o_1
XFILLER_0_78_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1627_ _0718_ VGND VGND VPWR VPWR _0772_ sky130_fd_sc_hd__buf_6
X_1558_ _0667_ VGND VGND VPWR VPWR _0673_ sky130_fd_sc_hd__buf_4
XTAP_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_354 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2530_ _1199_ net52 _0164_ _1211_ VGND VGND VPWR VPWR _0189_ sky130_fd_sc_hd__a211o_1
XFILLER_0_11_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2461_ _0836_ _1289_ _1462_ VGND VGND VPWR VPWR _0122_ sky130_fd_sc_hd__or3_1
XFILLER_0_51_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2392_ _1510_ _1528_ _1197_ VGND VGND VPWR VPWR _1529_ sky130_fd_sc_hd__o21ai_1
X_3013_ weights_inst.data_out\[13\] _0666_ VGND VGND VPWR VPWR _0671_ sky130_fd_sc_hd__and2_1
XFILLER_0_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2728_ _1244_ _0380_ _1125_ _0381_ _1342_ VGND VGND VPWR VPWR _0382_ sky130_fd_sc_hd__o311a_1
XFILLER_0_100_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2659_ _1345_ _1129_ _0209_ _0314_ _1287_ VGND VGND VPWR VPWR _0315_ sky130_fd_sc_hd__o311a_1
XFILLER_0_10_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1961_ _1036_ _1103_ VGND VGND VPWR VPWR _1104_ sky130_fd_sc_hd__nor2_1
XFILLER_0_83_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1892_ _0634_ VGND VGND VPWR VPWR _1036_ sky130_fd_sc_hd__buf_8
XFILLER_0_50_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2513_ _0716_ _0823_ _0790_ VGND VGND VPWR VPWR _0173_ sky130_fd_sc_hd__and3_1
XFILLER_0_51_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2444_ _0820_ _0829_ _1173_ VGND VGND VPWR VPWR _0105_ sky130_fd_sc_hd__and3_1
X_2375_ _1078_ _1392_ VGND VGND VPWR VPWR _1512_ sky130_fd_sc_hd__nor2_1
XFILLER_0_93_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_110 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2160_ net58 _0771_ VGND VGND VPWR VPWR _1301_ sky130_fd_sc_hd__nor2_2
X_2091_ _1232_ _0918_ _0851_ VGND VGND VPWR VPWR _1233_ sky130_fd_sc_hd__and3_1
XFILLER_0_88_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_cap1 _0653_ VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2993_ weights_inst.data_out\[3\] _0654_ _0658_ fsm_inst.done VGND VGND VPWR VPWR
+ net44 sky130_fd_sc_hd__a22o_1
XFILLER_0_61_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1944_ _1083_ _0856_ _1085_ _1086_ VGND VGND VPWR VPWR _1087_ sky130_fd_sc_hd__a31o_1
XFILLER_0_83_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1875_ _0713_ VGND VGND VPWR VPWR _1019_ sky130_fd_sc_hd__buf_4
XFILLER_0_9_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2427_ _0810_ _1439_ _1443_ VGND VGND VPWR VPWR _0089_ sky130_fd_sc_hd__or3_1
XFILLER_0_86_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2358_ _1298_ _1484_ _1486_ _1494_ _1396_ VGND VGND VPWR VPWR _1495_ sky130_fd_sc_hd__o311a_1
X_2289_ _0673_ _1416_ _1420_ _1427_ _0861_ VGND VGND VPWR VPWR _1428_ sky130_fd_sc_hd__o311a_1
XFILLER_0_94_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_308 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1660_ _0804_ VGND VGND VPWR VPWR _0805_ sky130_fd_sc_hd__clkbuf_8
X_1591_ net2 net3 VGND VGND VPWR VPWR _0736_ sky130_fd_sc_hd__and2b_1
XFILLER_0_40_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2212_ _0734_ _1146_ _1350_ _1351_ _1178_ VGND VGND VPWR VPWR _1352_ sky130_fd_sc_hd__a311o_1
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2143_ _1283_ _0725_ _1055_ VGND VGND VPWR VPWR _1284_ sky130_fd_sc_hd__or3b_1
XFILLER_0_56_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2074_ _1041_ _1213_ _1214_ _1215_ _0910_ VGND VGND VPWR VPWR _1216_ sky130_fd_sc_hd__a221o_1
XFILLER_0_88_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2976_ _1310_ _0640_ _0643_ _0952_ VGND VGND VPWR VPWR _0644_ sky130_fd_sc_hd__a211o_1
XFILLER_0_29_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1927_ _0952_ _1048_ _1058_ _1070_ VGND VGND VPWR VPWR _1071_ sky130_fd_sc_hd__o31a_1
X_1858_ _1000_ _1001_ VGND VGND VPWR VPWR _1002_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1789_ _0777_ VGND VGND VPWR VPWR _0934_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_99_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2830_ _0752_ _1182_ _0486_ _0487_ _1342_ VGND VGND VPWR VPWR _0488_ sky130_fd_sc_hd__o311a_1
XFILLER_0_58_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2761_ _1322_ _0388_ _0401_ _0414_ _0859_ VGND VGND VPWR VPWR _0012_ sky130_fd_sc_hd__o311a_1
XFILLER_0_26_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1712_ _0808_ _0856_ _0849_ VGND VGND VPWR VPWR _0857_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_5_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2692_ _1299_ _1302_ _1417_ _0346_ _0779_ VGND VGND VPWR VPWR _0347_ sky130_fd_sc_hd__o311a_1
XFILLER_0_53_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1643_ _0772_ _0787_ VGND VGND VPWR VPWR _0788_ sky130_fd_sc_hd__nor2_8
XANTENNA_1 _0137_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1574_ net3 _0718_ VGND VGND VPWR VPWR _0719_ sky130_fd_sc_hd__nand2b_4
XTAP_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2126_ _1117_ _0916_ VGND VGND VPWR VPWR _1267_ sky130_fd_sc_hd__nor2_1
X_2057_ _1041_ VGND VGND VPWR VPWR _1199_ sky130_fd_sc_hd__buf_4
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2959_ _1182_ _1224_ _1244_ VGND VGND VPWR VPWR _0626_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_17_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2813_ _1348_ _1516_ _0467_ _0468_ _1285_ VGND VGND VPWR VPWR _0469_ sky130_fd_sc_hd__o311a_1
XFILLER_0_81_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2744_ _1229_ _1399_ _1259_ VGND VGND VPWR VPWR _0398_ sky130_fd_sc_hd__a21o_1
XFILLER_0_14_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2675_ _0926_ _0713_ _0892_ VGND VGND VPWR VPWR _0331_ sky130_fd_sc_hd__and3_1
XFILLER_0_78_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1626_ _0765_ VGND VGND VPWR VPWR _0771_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_78_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1557_ _0661_ VGND VGND VPWR VPWR _0667_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_94_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2109_ _0915_ VGND VGND VPWR VPWR _1250_ sky130_fd_sc_hd__clkbuf_4
XTAP_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3089_ _0709_ VGND VGND VPWR VPWR _0055_ sky130_fd_sc_hd__inv_2
XFILLER_0_92_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_366 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2460_ _1365_ _0102_ _0108_ _0120_ VGND VGND VPWR VPWR _0121_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_51_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2391_ _1298_ _1514_ _1518_ _1527_ _0861_ VGND VGND VPWR VPWR _1528_ sky130_fd_sc_hd__o311a_1
XFILLER_0_48_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3012_ _0670_ VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__buf_1
XFILLER_0_74_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2727_ _1438_ _0221_ _1244_ VGND VGND VPWR VPWR _0381_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_73_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2658_ _0720_ _0901_ _1314_ _1256_ VGND VGND VPWR VPWR _0314_ sky130_fd_sc_hd__o31ai_1
X_2589_ _0800_ _1119_ _1467_ VGND VGND VPWR VPWR _0247_ sky130_fd_sc_hd__or3_1
XFILLER_0_10_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1609_ _0723_ VGND VGND VPWR VPWR _0754_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_69_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1960_ _0852_ _0785_ _0823_ VGND VGND VPWR VPWR _1103_ sky130_fd_sc_hd__and3_2
XFILLER_0_55_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1891_ _0915_ _1021_ _1024_ _1034_ VGND VGND VPWR VPWR _1035_ sky130_fd_sc_hd__a31o_1
XFILLER_0_43_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_391 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2512_ _1089_ _0790_ VGND VGND VPWR VPWR _0172_ sky130_fd_sc_hd__nand2_2
XFILLER_0_11_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2443_ _1343_ _0973_ _0912_ _1335_ VGND VGND VPWR VPWR _0104_ sky130_fd_sc_hd__a211o_1
X_2374_ _1117_ net52 VGND VGND VPWR VPWR _1511_ sky130_fd_sc_hd__and2_1
XFILLER_0_93_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_136 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_475 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_188 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2090_ _0825_ VGND VGND VPWR VPWR _1232_ sky130_fd_sc_hd__buf_4
XFILLER_0_45_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2992_ weights_inst.data_out\[2\] _0654_ _0658_ fsm_inst.done VGND VGND VPWR VPWR
+ net42 sky130_fd_sc_hd__a22o_1
XFILLER_0_90_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1943_ _0797_ _1084_ _0997_ _0754_ VGND VGND VPWR VPWR _1086_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_61_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1874_ _0915_ _1010_ _1017_ _0993_ VGND VGND VPWR VPWR _1018_ sky130_fd_sc_hd__a31o_1
XFILLER_0_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2426_ _1235_ _0962_ _1097_ VGND VGND VPWR VPWR _0088_ sky130_fd_sc_hd__or3b_1
XFILLER_0_86_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2357_ _1308_ _1488_ _1489_ _1493_ _1318_ VGND VGND VPWR VPWR _1494_ sky130_fd_sc_hd__a311o_4
XFILLER_0_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2288_ _0783_ _1421_ _1423_ _1426_ VGND VGND VPWR VPWR _1427_ sky130_fd_sc_hd__a31o_1
XFILLER_0_19_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1590_ _0711_ VGND VGND VPWR VPWR _0735_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_21_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2211_ _1199_ _1088_ _0879_ _0882_ _0725_ VGND VGND VPWR VPWR _1351_ sky130_fd_sc_hd__o2111a_1
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2142_ _0805_ _1275_ VGND VGND VPWR VPWR _1283_ sky130_fd_sc_hd__nor2_1
XFILLER_0_56_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2073_ net54 _0868_ VGND VGND VPWR VPWR _1215_ sky130_fd_sc_hd__nor2_1
XFILLER_0_72_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2975_ _0807_ _0641_ _0642_ _0778_ VGND VGND VPWR VPWR _0643_ sky130_fd_sc_hd__o211a_1
XFILLER_0_29_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1926_ _0782_ _1061_ _1062_ _1069_ _0993_ VGND VGND VPWR VPWR _1070_ sky130_fd_sc_hd__a311o_1
XFILLER_0_4_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1857_ _0826_ _0996_ VGND VGND VPWR VPWR _1001_ sky130_fd_sc_hd__nand2_4
XFILLER_0_44_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1788_ _0923_ _0925_ _0928_ _0932_ _0839_ VGND VGND VPWR VPWR _0933_ sky130_fd_sc_hd__o311a_1
X_2409_ _1113_ _1072_ _1150_ _1028_ VGND VGND VPWR VPWR _0071_ sky130_fd_sc_hd__a211o_1
XFILLER_0_98_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2760_ _0861_ _0402_ _1520_ _0413_ _0849_ VGND VGND VPWR VPWR _0414_ sky130_fd_sc_hd__a311o_1
XFILLER_0_53_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1711_ _0851_ _0855_ VGND VGND VPWR VPWR _0856_ sky130_fd_sc_hd__nand2_2
X_2691_ _0873_ _0344_ _0345_ VGND VGND VPWR VPWR _0346_ sky130_fd_sc_hd__or3_1
XFILLER_0_53_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1642_ _0729_ _0735_ VGND VGND VPWR VPWR _0787_ sky130_fd_sc_hd__nor2_8
XANTENNA_2 _0137_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1573_ _0717_ VGND VGND VPWR VPWR _0718_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_67_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2125_ _1123_ _0819_ _0975_ VGND VGND VPWR VPWR _1266_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_76_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2056_ _0934_ VGND VGND VPWR VPWR _1198_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_16_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2958_ _0578_ _0624_ _0843_ VGND VGND VPWR VPWR _0625_ sky130_fd_sc_hd__a21o_1
X_1909_ _0757_ _1052_ VGND VGND VPWR VPWR _1053_ sky130_fd_sc_hd__nor2_2
XFILLER_0_44_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2889_ _0801_ _0890_ _1150_ _0550_ _0782_ VGND VGND VPWR VPWR _0551_ sky130_fd_sc_hd__o311a_1
XFILLER_0_32_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput50 net50 VGND VGND VPWR VPWR wbs_dat_o[9] sky130_fd_sc_hd__buf_12
XFILLER_0_37_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2812_ _0936_ _0888_ _0124_ VGND VGND VPWR VPWR _0468_ sky130_fd_sc_hd__or3_1
XFILLER_0_26_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2743_ _1190_ _0214_ _1244_ VGND VGND VPWR VPWR _0397_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_14_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2674_ _1274_ _0871_ _0181_ VGND VGND VPWR VPWR _0330_ sky130_fd_sc_hd__nand3_1
XFILLER_0_78_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1625_ _0769_ VGND VGND VPWR VPWR _0770_ sky130_fd_sc_hd__buf_6
XFILLER_0_41_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1556_ _0516_ _0580_ VGND VGND VPWR VPWR _0661_ sky130_fd_sc_hd__xor2_4
XFILLER_0_94_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2108_ _1204_ _0758_ VGND VGND VPWR VPWR _1249_ sky130_fd_sc_hd__nor2_4
XTAP_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3088_ _0709_ VGND VGND VPWR VPWR _0054_ sky130_fd_sc_hd__inv_2
X_2039_ _0772_ _0946_ VGND VGND VPWR VPWR _1181_ sky130_fd_sc_hd__nor2_4
XFILLER_0_92_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2390_ _1310_ _1521_ _1522_ _1526_ _1318_ VGND VGND VPWR VPWR _1527_ sky130_fd_sc_hd__a311o_1
X_3011_ weights_inst.data_out\[12\] _0666_ VGND VGND VPWR VPWR _0670_ sky130_fd_sc_hd__and2_1
XFILLER_0_58_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2726_ _0771_ _0896_ VGND VGND VPWR VPWR _0380_ sky130_fd_sc_hd__nor2_2
XFILLER_0_6_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2657_ _0655_ _0989_ VGND VGND VPWR VPWR _0313_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1608_ _0722_ _0734_ _0748_ _0752_ VGND VGND VPWR VPWR _0753_ sky130_fd_sc_hd__a22o_1
X_2588_ _0751_ _1294_ _1500_ _0245_ _1047_ VGND VGND VPWR VPWR _0246_ sky130_fd_sc_hd__o311a_1
X_1539_ net6 net8 VGND VGND VPWR VPWR _0484_ sky130_fd_sc_hd__nand2_1
XTAP_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1890_ _0694_ _1029_ _1033_ _0841_ VGND VGND VPWR VPWR _1034_ sky130_fd_sc_hd__a31o_1
XFILLER_0_3_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2511_ _0836_ _1315_ _1277_ VGND VGND VPWR VPWR _0171_ sky130_fd_sc_hd__or3_4
XFILLER_0_11_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2442_ _1089_ _1343_ _0929_ _0942_ VGND VGND VPWR VPWR _0103_ sky130_fd_sc_hd__a31o_1
X_2373_ _1273_ _1499_ _1503_ _1509_ _1396_ VGND VGND VPWR VPWR _1510_ sky130_fd_sc_hd__o311a_1
XFILLER_0_75_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2709_ _1356_ _0360_ _0363_ _0860_ VGND VGND VPWR VPWR _0364_ sky130_fd_sc_hd__a211o_1
XFILLER_0_100_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_395 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2991_ weights_inst.data_out\[1\] _0654_ net53 fsm_inst.batch_norm_en VGND VGND VPWR
+ VPWR net31 sky130_fd_sc_hd__a22o_1
XFILLER_0_28_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1942_ _0819_ _1084_ VGND VGND VPWR VPWR _1085_ sky130_fd_sc_hd__nand2_1
XFILLER_0_83_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1873_ _1011_ _1014_ _1016_ _0890_ _0922_ VGND VGND VPWR VPWR _1017_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_43_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2425_ _1165_ _0085_ _0086_ _0744_ _0839_ VGND VGND VPWR VPWR _0087_ sky130_fd_sc_hd__o221a_1
X_2356_ _0945_ _1002_ _1490_ _1492_ _0978_ VGND VGND VPWR VPWR _1493_ sky130_fd_sc_hd__o311a_1
X_2287_ _1047_ _1424_ _1425_ _0842_ VGND VGND VPWR VPWR _1426_ sky130_fd_sc_hd__a31o_1
XFILLER_0_29_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2210_ _1136_ _1173_ VGND VGND VPWR VPWR _1350_ sky130_fd_sc_hd__nand2_2
X_2141_ _1232_ _0770_ _0854_ VGND VGND VPWR VPWR _1282_ sky130_fd_sc_hd__and3_1
X_2072_ _0784_ _0743_ _0903_ VGND VGND VPWR VPWR _1214_ sky130_fd_sc_hd__or3_2
XFILLER_0_88_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2974_ _1013_ _1314_ _0303_ _0985_ VGND VGND VPWR VPWR _0642_ sky130_fd_sc_hd__a211o_1
XFILLER_0_29_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1925_ _1063_ _0722_ _1065_ _1068_ _0914_ VGND VGND VPWR VPWR _1069_ sky130_fd_sc_hd__a311oi_4
XFILLER_0_56_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1856_ _0999_ VGND VGND VPWR VPWR _1000_ sky130_fd_sc_hd__buf_4
X_1787_ _0788_ _0929_ _0931_ _0836_ VGND VGND VPWR VPWR _0932_ sky130_fd_sc_hd__a211o_1
XFILLER_0_4_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2408_ _1110_ _1020_ _0911_ VGND VGND VPWR VPWR _0070_ sky130_fd_sc_hd__a21o_1
X_2339_ _0914_ _1474_ _1476_ _0661_ VGND VGND VPWR VPWR _1477_ sky130_fd_sc_hd__a31o_1
XFILLER_0_67_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2690_ _0939_ _0831_ _0897_ VGND VGND VPWR VPWR _0345_ sky130_fd_sc_hd__and3_2
X_1710_ _0852_ _0740_ _0854_ VGND VGND VPWR VPWR _0855_ sky130_fd_sc_hd__and3_4
X_1641_ _0785_ VGND VGND VPWR VPWR _0786_ sky130_fd_sc_hd__buf_4
XANTENNA_3 _0177_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1572_ net2 VGND VGND VPWR VPWR _0717_ sky130_fd_sc_hd__clkbuf_8
XTAP_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2124_ _0718_ _0727_ _0946_ VGND VGND VPWR VPWR _1265_ sky130_fd_sc_hd__and3_4
XFILLER_0_83_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2055_ _0848_ VGND VGND VPWR VPWR _1197_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_16_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_251 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2957_ _0579_ _0622_ _0703_ VGND VGND VPWR VPWR _0624_ sky130_fd_sc_hd__a21o_1
XFILLER_0_32_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2888_ _1019_ _1043_ _1206_ _0172_ _1140_ VGND VGND VPWR VPWR _0550_ sky130_fd_sc_hd__a221o_1
X_1908_ _0765_ _0831_ VGND VGND VPWR VPWR _1052_ sky130_fd_sc_hd__nor2_2
XFILLER_0_44_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1839_ _0959_ VGND VGND VPWR VPWR _0983_ sky130_fd_sc_hd__buf_4
XFILLER_0_32_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput40 net40 VGND VGND VPWR VPWR wbs_dat_o[28] sky130_fd_sc_hd__buf_12
XFILLER_0_53_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2811_ _0769_ _0999_ _0851_ VGND VGND VPWR VPWR _0467_ sky130_fd_sc_hd__and3_2
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2742_ _1244_ _1072_ _0109_ _0395_ _0783_ VGND VGND VPWR VPWR _0396_ sky130_fd_sc_hd__o311a_1
XFILLER_0_26_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2673_ _0873_ _0747_ _1065_ VGND VGND VPWR VPWR _0329_ sky130_fd_sc_hd__or3b_1
X_1624_ _0768_ VGND VGND VPWR VPWR _0769_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_78_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1555_ _0645_ VGND VGND VPWR VPWR _0655_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_94_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3087_ _0709_ VGND VGND VPWR VPWR _0053_ sky130_fd_sc_hd__inv_2
X_2107_ _0810_ _1247_ VGND VGND VPWR VPWR _1248_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2038_ _0750_ VGND VGND VPWR VPWR _1180_ sky130_fd_sc_hd__buf_4
XFILLER_0_76_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3010_ _0669_ VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__buf_1
XFILLER_0_78_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_308 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2725_ _0752_ _0377_ _0378_ _0783_ VGND VGND VPWR VPWR _0379_ sky130_fd_sc_hd__o211a_1
XFILLER_0_42_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2656_ _0306_ _0311_ _1365_ VGND VGND VPWR VPWR _0312_ sky130_fd_sc_hd__a21oi_1
X_1607_ _0751_ VGND VGND VPWR VPWR _0752_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2587_ _0878_ _0713_ _0971_ _1166_ _1060_ VGND VGND VPWR VPWR _0245_ sky130_fd_sc_hd__a311o_1
XFILLER_0_59_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1538_ net6 net4 net58 _0462_ VGND VGND VPWR VPWR _0473_ sky130_fd_sc_hd__a31o_4
XTAP_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_500 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2510_ _0810_ _0940_ _1084_ VGND VGND VPWR VPWR _0170_ sky130_fd_sc_hd__or3_1
XFILLER_0_3_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2441_ _0706_ _0099_ _0101_ _1164_ VGND VGND VPWR VPWR _0102_ sky130_fd_sc_hd__a211o_1
XFILLER_0_59_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2372_ _0779_ _1504_ _1505_ _1508_ _0667_ VGND VGND VPWR VPWR _1509_ sky130_fd_sc_hd__a311o_1
XFILLER_0_91_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2708_ _0963_ _0361_ _0362_ VGND VGND VPWR VPWR _0363_ sky130_fd_sc_hd__and3_1
XFILLER_0_100_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2639_ _1109_ _1236_ _1523_ _0295_ _0782_ VGND VGND VPWR VPWR _0296_ sky130_fd_sc_hd__o311a_1
XFILLER_0_100_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2990_ weights_inst.data_out\[0\] _0654_ net53 fsm_inst.cnn_en VGND VGND VPWR VPWR
+ net20 sky130_fd_sc_hd__a22o_1
XFILLER_0_28_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1941_ _0784_ _0868_ VGND VGND VPWR VPWR _1084_ sky130_fd_sc_hd__nor2_4
XFILLER_0_61_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1872_ _0741_ _1015_ VGND VGND VPWR VPWR _1016_ sky130_fd_sc_hd__nor2_4
XFILLER_0_56_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_138 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2424_ _1011_ _0971_ _0973_ _0750_ VGND VGND VPWR VPWR _0086_ sky130_fd_sc_hd__a31o_1
XFILLER_0_86_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2355_ _1000_ _1043_ _1491_ _0800_ VGND VGND VPWR VPWR _1492_ sky130_fd_sc_hd__a211o_1
X_2286_ _0947_ _0948_ _1314_ _1083_ VGND VGND VPWR VPWR _1425_ sky130_fd_sc_hd__a211o_1
XFILLER_0_79_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_116 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2140_ _1109_ VGND VGND VPWR VPWR _1281_ sky130_fd_sc_hd__buf_4
X_2071_ _0887_ _0959_ VGND VGND VPWR VPWR _1213_ sky130_fd_sc_hd__and2_4
XFILLER_0_88_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_327 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2973_ _1211_ _1120_ VGND VGND VPWR VPWR _0641_ sky130_fd_sc_hd__nand2_1
X_1924_ _1066_ _0864_ _1067_ VGND VGND VPWR VPWR _1068_ sky130_fd_sc_hd__and3b_1
XFILLER_0_17_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1855_ _0998_ VGND VGND VPWR VPWR _0999_ sky130_fd_sc_hd__buf_4
XFILLER_0_24_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1786_ _0727_ _0930_ VGND VGND VPWR VPWR _0931_ sky130_fd_sc_hd__nor2_8
XFILLER_0_12_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2407_ _1391_ _0880_ _0900_ VGND VGND VPWR VPWR _0069_ sky130_fd_sc_hd__or3_1
XFILLER_0_99_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2338_ _0799_ _1475_ _1054_ VGND VGND VPWR VPWR _1476_ sky130_fd_sc_hd__or3b_1
X_2269_ _1367_ _1025_ _1407_ _1040_ VGND VGND VPWR VPWR _1408_ sky130_fd_sc_hd__a211o_1
XFILLER_0_46_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1640_ _0784_ VGND VGND VPWR VPWR _0785_ sky130_fd_sc_hd__clkbuf_8
XANTENNA_4 _0204_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1571_ _0715_ VGND VGND VPWR VPWR _0716_ sky130_fd_sc_hd__buf_4
XFILLER_0_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2123_ _0985_ VGND VGND VPWR VPWR _1264_ sky130_fd_sc_hd__buf_4
XFILLER_0_88_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2054_ _1160_ _1163_ _1195_ _0861_ VGND VGND VPWR VPWR _1196_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_49_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2956_ _0744_ _1130_ _1261_ VGND VGND VPWR VPWR _0622_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_29_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2887_ _0923_ _0546_ _0547_ _1047_ VGND VGND VPWR VPWR _0549_ sky130_fd_sc_hd__o211a_1
X_1907_ _1049_ _0979_ _1050_ VGND VGND VPWR VPWR _1051_ sky130_fd_sc_hd__or3_1
XFILLER_0_44_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1838_ _0751_ _0974_ _0977_ _0978_ _0981_ VGND VGND VPWR VPWR _0982_ sky130_fd_sc_hd__o311a_1
XFILLER_0_4_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1769_ _0776_ VGND VGND VPWR VPWR _0914_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_12_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput30 net30 VGND VGND VPWR VPWR wbs_dat_o[19] sky130_fd_sc_hd__buf_12
Xoutput41 net41 VGND VGND VPWR VPWR wbs_dat_o[29] sky130_fd_sc_hd__buf_12
XFILLER_0_101_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2810_ _1298_ _0463_ _0465_ _1039_ VGND VGND VPWR VPWR _0466_ sky130_fd_sc_hd__o31a_1
XFILLER_0_54_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2741_ _1124_ _1229_ _1072_ _0803_ _1261_ VGND VGND VPWR VPWR _0395_ sky130_fd_sc_hd__a221o_1
XFILLER_0_81_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2672_ _1403_ _1088_ _1027_ _0327_ _1285_ VGND VGND VPWR VPWR _0328_ sky130_fd_sc_hd__o311a_1
XFILLER_0_10_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1623_ _0715_ VGND VGND VPWR VPWR _0768_ sky130_fd_sc_hd__buf_4
XFILLER_0_22_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1554_ _0634_ VGND VGND VPWR VPWR _0645_ sky130_fd_sc_hd__buf_6
.ends

